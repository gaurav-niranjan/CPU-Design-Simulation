//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "try.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w58;    //: /sn:0 {0}(-133,-414)(-133,-505){1}
reg [7:0] w65;    //: /sn:0 {0}(#:-301,-458)(-272,-458)(-272,-511){1}
reg w50;    //: /sn:0 {0}(-662,-188)(-559,-188)(-559,-208)(-540,-208){1}
reg w71;    //: /sn:0 {0}(6,-37)(6,-39)(101,-39)(101,-67)(114,-67)(114,-49)(129,-49)(129,-59){1}
reg w19;    //: /sn:0 {0}(673,446)(646,446)(646,443)(636,443){1}
reg w66;    //: /sn:0 {0}(775,-382)(775,-422)(774,-422)(774,-437){1}
//: {2}(776,-439)(803,-439){3}
//: {4}(774,-441)(774,-461)(712,-461)(712,-480){5}
reg w73;    //: /sn:0 {0}(-42,104)(-42,94)(-1,94)(-1,13){1}
reg w63;    //: /sn:0 {0}(705,-547)(705,-542){1}
//: {2}(703,-540)(695,-540)(695,-580){3}
//: {4}(705,-538)(705,-530){5}
reg w52;    //: /sn:0 {0}(-126,-572)(-126,-567){1}
//: {2}(-128,-565)(-143,-565)(-143,-587){3}
//: {4}(-126,-563)(-126,-555){5}
reg w17;    //: /sn:0 {0}(337,457)(337,467)(307,467)(307,472){1}
reg w67;    //: /sn:0 {0}(697,-399)(697,-470)(698,-470)(698,-480){1}
reg w14;    //: /sn:0 {0}(-600,-228)(-540,-228){1}
reg w69;    //: /sn:0 {0}(82,112)(82,72)(115,72)(115,-5){1}
//: {2}(117,-7)(144,-7){3}
//: {4}(113,-7)(81,-7)(81,34)(13,34)(13,13){5}
reg w78;    //: /sn:0 {0}(1414,-168)(1414,-272)(1352,-272)(1352,-291){1}
reg w15;    //: /sn:0 {0}(372,229)(394,229)(394,221){1}
reg [7:0] w5;    //: /sn:0 {0}(#:165,483)(278,483)(278,480)(293,480){1}
reg w61;    //: /sn:0 {0}(-280,-525)(-329,-525)(-329,-526)(-344,-526){1}
reg w43;    //: /sn:0 {0}(-510,25)(-431,25)(-431,39)(-416,39){1}
reg w76;    //: /sn:0 {0}(1338,-190)(1338,-182)(1339,-182)(1339,-134){1}
reg w40;    //: /sn:0 {0}(-593,-12)(-653,-12)(-653,-132)(-662,-132){1}
reg w57;    //: /sn:0 {0}(-57,-403)(-57,-462){1}
//: {2}(-55,-464)(-28,-464){3}
//: {4}(-57,-466)(-57,-486)(-119,-486)(-119,-505){5}
reg w77;    //: /sn:0 {0}(1345,-341)(1345,-370){1}
//: {2}(1347,-372)(1530,-372){3}
//: {4}(1345,-374)(1345,-398)(1333,-398)(1333,-413){5}
wire w6;    //: /sn:0 {0}(907,53)(907,80)(859,80){1}
wire w13;    //: /sn:0 {0}(545,-25)(477,-25)(477,179){1}
//: {2}(479,181)(798,181){3}
//: {4}(477,183)(477,193)(410,193){5}
wire w16;    //: /sn:0 {0}(545,47)(509,47)(509,138){1}
//: {2}(511,140)(798,140){3}
//: {4}(509,142)(509,204)(410,204){5}
wire w7;    //: /sn:0 {0}(753,402)(640,402)(640,343)(562,343){1}
wire [2:0] w34;    //: /sn:0 {0}(293,512)(258,512)(#:258,441)(#:224,441){1}
wire w59;    //: /sn:0 {0}(-12,-464)(51,-464)(51,-451){1}
wire w25;    //: /sn:0 {0}(912,53)(912,84)(905,84)(905,98){1}
wire w39;    //: /sn:0 {0}(-502,-105)(-549,-105)(-549,10){1}
wire [3:0] w4;    //: /sn:0 {0}(#:110,208)(264,208){1}
//: {2}(268,208)(#:273,208)(273,199)(381,199){3}
//: {4}(266,206)(266,194){5}
wire [7:0] w62;    //: /sn:0 {0}(874,-421)(842,-421)(#:842,-497)(753,-497)(753,-507)(#:722,-507){1}
wire [7:0] w72;    //: /sn:0 {0}(212,52)(51,52)(51,-14)(#:23,-14){1}
wire w56;    //: /sn:0 {0}(-371,410)(-300,410){1}
//: {2}(-296,410)(423,410)(423,225)(410,225){3}
//: {4}(-298,408)(-298,370){5}
wire [7:0] w36;    //: /sn:0 {0}(#:1150,-36)(1181,-36)(1181,42)(#:1606,42)(1606,-216){1}
//: {2}(1608,-218)(#:1661,-218){3}
//: {4}(1606,-220)(1606,-308)(1582,-308){5}
wire w82;    //: /sn:0 {0}(410,186)(453,186)(453,127){1}
//: {2}(455,125)(798,125){3}
//: {4}(453,123)(453,-61)(545,-61){5}
wire [2:0] w0;    //: /sn:0 {0}(#:110,309)(184,309){1}
//: {2}(188,309)(301,309)(301,310){3}
//: {4}(303,312)(440,312){5}
//: {6}(301,314)(301,330){7}
//: {8}(#:186,311)(186,441)(208,441){9}
wire w3;    //: /sn:0 {0}(110,269)(211,269){1}
//: {2}(215,269)(311,269){3}
//: {4}(315,269)(337,269){5}
//: {6}(313,271)(313,296)(366,296){7}
//: {8}(213,271)(213,305)(216,305)(216,436){9}
wire w22;    //: /sn:0 {0}(410,214)(422,214)(422,-169)(-174,-169)(-174,-164){1}
//: {2}(-176,-162)(-545,-162)(-545,-154)(-632,-154)(-632,16){3}
//: {4}(-174,-160)(-174,-137)(-221,-137){5}
wire w20;    //: /sn:0 {0}(-371,426)(-322,426){1}
//: {2}(-318,426)(429,426)(429,221)(410,221){3}
//: {4}(-320,424)(-320,382)(-319,382)(-319,371){5}
wire [7:0] w60;    //: /sn:0 {0}(#:1362,-318)(1393,-318)(1393,-308)(#:1566,-308){1}
wire w29;    //: /sn:0 {0}(753,311)(613,311)(613,316)(562,316){1}
wire w30;    //: /sn:0 {0}(753,282)(694,282)(694,297)(665,297)(665,309)(562,309){1}
wire w42;    //: /sn:0 {0}(348,524)(307,524)(307,520){1}
wire [7:0] w37;    //: /sn:0 {0}(#:545,-107)(-140,-107){1}
//: {2}(-144,-107)(-181,-107)(-181,-106)(-195,-106){3}
//: {4}(-199,-106)(-209,-106)(-209,-105)(-221,-105){5}
//: {6}(-197,-104)(#:-197,-94)(-198,-94)(-198,-80){7}
//: {8}(-142,-105)(-142,-49){9}
//: {10}(-144,-47)(-164,-47){11}
//: {12}(-142,-45)(#:-142,550)(483,550){13}
//: {14}(487,550)(510,550)(510,548)(522,548){15}
//: {16}(526,548)(563,548){17}
//: {18}(524,550)(#:524,560)(525,560)(525,617){19}
//: {20}(485,548)(#:485,532){21}
wire [7:0] w18;    //: /sn:0 {0}(#:322,496)(357,496)(357,441)(475,441)(#:475,503){1}
wire w12;    //: /sn:0 {0}(545,-43)(466,-43)(466,128){1}
//: {2}(468,130)(798,130){3}
//: {4}(466,132)(466,190)(410,190){5}
wire [7:0] w10;    //: /sn:0 {0}(#:6,354)(106,354)(106,309){1}
//: {2}(106,308)(106,269){3}
//: {4}(106,268)(106,208){5}
//: {6}(106,207)(106,162)(362,162)(362,116)(#:347,116)(347,58)(335,58)(335,52)(#:228,52){7}
wire w23;    //: /sn:0 {0}(382,296)(410,296){1}
//: {2}(414,296)(448,296)(448,307){3}
//: {4}(412,298)(412,504){5}
//: {6}(410,506)(400,506)(400,507)(385,507){7}
//: {8}(412,508)(412,519)(462,519){9}
wire w91;    //: /sn:0 {0}(545,-85)(435,-85)(435,118){1}
//: {2}(437,120)(798,120){3}
//: {4}(435,122)(435,179)(410,179){5}
wire w54;    //: /sn:0 {0}(819,168)(871,168)(871,150)(886,150){1}
wire w70;    //: /sn:0 {0}(160,-7)(220,-7)(220,47){1}
wire w84;    //: /sn:0 {0}(-577,-12)(-494,-12)(-494,15)(-510,15){1}
wire [7:0] w86;    //: /sn:0 {0}(495,503)(495,468)(#:1187,468)(1187,340){1}
//: {2}(1189,338)(#:1199,338)(1199,339)(1222,339){3}
//: {4}(1187,336)(1187,237){5}
//: {6}(1187,233)(1187,225){7}
//: {8}(1185,235)(#:1177,235)(1177,212)(1088,212){9}
wire w24;    //: /sn:0 {0}(917,53)(917,136)(939,136)(939,146){1}
//: {2}(941,148)(960,148){3}
//: {4}(964,148)(1134,148)(1134,460)(546,460)(546,342){5}
//: {6}(962,146)(962,-140)(1160,-140)(1160,-198)(1333,-198){7}
//: {8}(937,148)(907,148){9}
wire [7:0] w21;    //: /sn:0 {0}(-12,-12)(-74,-12)(#:-74,-55)(-126,-55)(#:-126,-233)(-37,-233)(-37,-249)(-65,-249){1}
//: {2}(-67,-251)(-67,-301)(-240,-301)(-240,-511){3}
//: {4}(-69,-249)(-132,-249){5}
//: {6}(-134,-251)(-134,-274){7}
//: {8}(-136,-249)(#:-181,-249){9}
wire [2:0] w1;    //: /sn:0 {0}(#:456,312)(498,312){1}
//: {2}(502,312)(522,312)(522,320)(533,320){3}
//: {4}(#:500,314)(500,422)(753,422){5}
wire w31;    //: /sn:0 {0}(753,260)(652,260)(652,274)(593,274)(593,303)(562,303){1}
wire w32;    //: /sn:0 {0}(562,296)(587,296)(587,266)(630,266)(630,240)(753,240){1}
wire w68;    //: /sn:0 {0}(819,-439)(882,-439)(882,-426){1}
wire [7:0] w53;    //: /sn:0 {0}(119,-389)(109,-389)(109,-404)(#:120,-404)(120,-444){1}
//: {2}(122,-446)(229,-446)(229,-467)(270,-467){3}
//: {4}(274,-467)(340,-467){5}
//: {6}(344,-467)(355,-467)(355,-316)(1327,-316){7}
//: {8}(#:342,-469)(342,-505)(687,-505){9}
//: {10}(272,-465)(#:272,-318)(-576,-318)(-576,-245)(-540,-245){11}
//: {12}(118,-446)(#:59,-446){13}
wire w8;    //: /sn:0 {0}(753,385)(645,385)(645,336)(562,336){1}
wire w46;    //: /sn:0 {0}(410,211)(530,211)(530,158){1}
//: {2}(532,156)(798,156){3}
//: {4}(530,154)(530,104)(545,104){5}
wire [7:0] w27;    //: /sn:0 {0}(#:579,548)(1091,548)(1091,-26)(1121,-26){1}
wire w44;    //: /sn:0 {0}(-624,21)(-603,21)(-603,20)(-586,20){1}
wire w75;    //: /sn:0 {0}(1338,-206)(1338,-291){1}
wire w35;    //: /sn:0 {0}(-371,378)(-357,378)(-357,347)(-549,347)(-549,114){1}
//: {2}(-547,112)(-537,112)(-537,113)(-513,113){3}
//: {4}(-549,110)(-549,31){5}
wire w28;    //: /sn:0 {0}(753,338)(717,338)(717,323)(562,323){1}
wire w80;    //: /sn:0 {0}(-754,426)(-765,426)(-765,348)(-729,348)(-729,-258)(-719,-258)(-719,-264)(-628,-264){1}
//: {2}(-624,-264)(-540,-264){3}
//: {4}(-626,-266)(-626,-324){5}
wire w49;    //: /sn:0 {0}(545,25)(498,25)(498,159){1}
//: {2}(500,161)(798,161){3}
//: {4}(498,163)(498,200)(410,200){5}
wire w45;    //: /sn:0 {0}(819,132)(871,132)(871,145)(886,145){1}
wire w11;    //: /sn:0 {0}(753,365)(689,365)(689,329)(562,329){1}
wire [7:0] w48;    //: /sn:0 {0}(#:784,-93)(1094,-93)(1094,-46)(1121,-46){1}
wire [7:0] w2;    //: /sn:0 {0}(#:628,216)(672,216){1}
//: {2}(676,216)(#:686,216)(686,211)(753,211){3}
//: {4}(674,214)(#:674,205){5}
wire w74;    //: /sn:0 {0}(1546,-372)(1559,-372)(1559,-293)(1574,-293)(1574,-303){1}
wire w41;    //: /sn:0 {0}(689,446)(725,446)(725,438)(753,438){1}
wire w47;    //: /sn:0 {0}(545,-1)(488,-1)(488,141){1}
//: {2}(490,143)(502,143)(502,135)(798,135){3}
//: {4}(488,145)(488,197)(410,197){5}
wire w83;    //: /sn:0 {0}(545,63)(518,63)(518,164){1}
//: {2}(520,166)(798,166){3}
//: {4}(518,168)(518,207)(410,207){5}
wire w94;    //: /sn:0 {0}(410,218)(426,218)(426,394)(-245,394){1}
//: {2}(-247,392)(-247,364){3}
//: {4}(-249,394)(-371,394){5}
wire w92;    //: /sn:0 {0}(410,176)(577,176)(577,173){1}
//: {2}(579,171)(753,171){3}
//: {4}(757,171)(798,171){5}
//: {6}(755,169)(755,80)(843,80){7}
//: {8}(575,171)(565,171)(565,186)(576,186)(576,488){9}
//: {10}(574,490)(558,490)(558,510)(548,510)(548,496){11}
//: {12}(576,492)(576,533)(571,533)(571,543){13}
wire [7:0] w38;    //: /sn:0 {0}(43,-446)(11,-446)(#:11,-522)(-78,-522)(-78,-532)(#:-109,-532){1}
wire [7:0] w55;    //: /sn:0 {0}(-144,-530)(-172,-530)(-172,-552)(-217,-552)(-217,-609)(#:-256,-609)(#:-256,-540){1}
wire w64;    //: /sn:0 {0}(-232,-525)(-212,-525)(-212,-512)(-190,-512){1}
wire w26;    //: /sn:0 {0}(912,32)(912,2)(1137,2)(1137,-13){1}
wire w9;    //: /sn:0 {0}(545,-73)(441,-73)(441,150){1}
//: {2}(443,152)(553,152)(553,145)(798,145){3}
//: {4}(441,154)(441,183)(410,183){5}
wire w93;    //: /sn:0 {0}(410,172)(553,172)(553,179)(693,179){1}
//: {2}(695,177)(695,176)(786,176){3}
//: {4}(790,176)(798,176){5}
//: {6}(788,174)(788,164)(913,164)(913,139)(905,139)(905,114){7}
//: {8}(695,181)(695,197)(691,197){9}
//: {10}(687,197)(679,197){11}
//: {12}(689,199)(689,206)(681,206)(681,441){13}
wire w79;    //: /sn:0 {0}(-669,50)(-669,21)(-640,21){1}
wire [7:0] w51;    //: /sn:0 {0}(#:890,-421)(900,-421)(900,-341)(602,-341)(602,-226)(666,-226)(666,-164){1}
//: {2}(#:668,-162)(681,-162)(681,-227)(718,-227){3}
//: {4}(666,-160)(666,-124){5}
//: {6}(#:668,-122)(674,-122)(674,189){7}
//: {8}(664,-122)(222,-122)(222,-121)(-221,-121){9}
//: {10}(666,-120)(666,-115)(535,-115)(535,-96)(#:545,-96){11}
//: enddecls

  //: comment g116 @(1239,-340) /sn:0 /R:14
  //: /line:"Address to write"
  //: /end
  _GGBUFIF3 #(4, 6) g8 (.Z(w1), .I(w0), .E(w23));   //: @(446,312) /sn:0 /w:[ 0 5 3 ]
  //: LED g4 (w4) @(266,187) /sn:0 /w:[ 5 ] /type:1
  _GGBUFIF3 #(4, 6) g17 (.Z(w34), .I(w0), .E(w3));   //: @(214,441) /sn:0 /w:[ 1 9 9 ]
  //: joint g137 (w93) @(788, 176) /w:[ 4 6 3 -1 ]
  //: joint g92 (w63) @(705, -540) /w:[ -1 1 2 4 ]
  _GGRAM8x8 #(10, 60, 70, 10, 10, 10) g74 (.A(w55), .D(w38), .WE(w52), .OE(w57), .CS(w58));   //: @(-126,-531) /w:[ 0 1 5 5 1 ]
  comparator g30 (.input_1(w37), .input_2(w51), .comparator_enable(w22), .comparator_result(w39));   //: @(-500, -153) /sz:(279, 64) /R:2 /sn:0 /p:[ Ri0>5 Ri1>9 Ri2>5 Lo0<0 ]
  //: SWITCH g130 (w19) @(619,443) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: frame g1 @(-89,-94) /sn:0 /wi:325 /ht:237 /tx:"RAM_READ"
  //: joint g77 (w57) @(-57, -464) /w:[ 2 4 -1 1 ]
  //: SWITCH g111 (w77) @(1333,-426) /sn:0 /R:3 /w:[ 5 ] /st:0 /dn:1
  _GGNBUF #(2) g144 (.I(w40), .Z(w84));   //: @(-587,-12) /sn:0 /w:[ 0 0 ]
  //: joint g51 (w12) @(466, 130) /w:[ 2 1 -1 4 ]
  //: LED g70 (w35) @(-506,113) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: joint g149 (w20) @(-320, 426) /w:[ 2 4 1 -1 ]
  //: joint g25 (w36) @(1606, -218) /w:[ 2 4 -1 1 ]
  _GGBUFIF #(4, 6) g103 (.Z(w75), .I(w76), .E(w24));   //: @(1338,-196) /sn:0 /R:1 /w:[ 0 0 7 ]
  //: comment g10 @(314,336) /sn:0
  //: /line:"Register/Immediate value"
  //: /line:""
  //: /end
  //: SWITCH g65 (w14) @(-617,-228) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g64 (w42) @(355,524) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: joint g72 (w80) @(-626, -264) /w:[ 2 4 1 -1 ]
  //: joint g49 (w9) @(441, 152) /w:[ 2 1 -1 4 ]
  //: comment g142 @(-751,-197) /sn:0
  //: /line:"PC_CLOCK"
  //: /end
  _GGNBUF #(2) g136 (.I(w93), .Z(w25));   //: @(905,108) /sn:0 /R:1 /w:[ 7 1 ]
  //: joint g6 (w4) @(266, 208) /w:[ 2 4 1 -1 ]
  //: LED g7 (w3) @(344,269) /sn:0 /R:3 /w:[ 5 ] /type:1
  _GGCLOCK_P100_0_50 g35 (.Z(w79));   //: @(-669,65) /sn:0 /R:1 /w:[ 0 ] /omega:100 /phi:0 /duty:50
  _GGOR2 #(6) g58 (.I0(w45), .I1(w54), .Z(w24));   //: @(897,148) /sn:0 /w:[ 1 1 9 ]
  //: joint g56 (w83) @(518, 166) /w:[ 2 1 -1 4 ]
  //: LED g124 (w37) @(-171,-47) /sn:0 /R:1 /w:[ 11 ] /type:1
  //: SWITCH g98 (w69) @(82,126) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g85 (w61) @(-361,-526) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: LED g67 (w21) @(-134,-281) /sn:0 /w:[ 7 ] /type:1
  //: LED g126 (w37) @(-198,-73) /sn:0 /R:2 /w:[ 7 ] /type:1
  //: SWITCH g33 (w43) @(-398,39) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  //: joint g54 (w49) @(498, 161) /w:[ 2 1 -1 4 ]
  //: SWITCH g81 (w52) @(-143,-600) /sn:0 /R:3 /w:[ 3 ] /st:1 /dn:1
  _GGBUFIF8 #(4, 6) g40 (.Z(w2), .I(w51), .E(w93));   //: @(674,195) /sn:0 /R:3 /w:[ 5 7 11 ]
  //: joint g52 (w13) @(477, 181) /w:[ 2 1 -1 4 ]
  //: joint g132 (w86) @(1187, 338) /w:[ 2 4 -1 1 ]
  _GGBUFIF #(4, 6) g108 (.Z(w41), .I(w19), .E(w93));   //: @(679,446) /sn:0 /w:[ 0 0 13 ]
  //: joint g12 (w3) @(313, 269) /w:[ 4 -1 3 6 ]
  //: LED g131 (w86) @(1229,339) /sn:0 /R:3 /w:[ 3 ] /type:1
  _GGRAM8x8 #(10, 60, 70, 10, 10, 10) g106 (.A(w53), .D(w60), .WE(w77), .OE(w78), .CS(w75));   //: @(1345,-317) /w:[ 7 0 0 1 1 ]
  _GGRAM8x8 #(10, 60, 70, 10, 10, 10) g96 (.A(w21), .D(w72), .WE(w71), .OE(w69), .CS(w73));   //: @(6,-13) /w:[ 0 1 0 5 1 ]
  //: comment g117 @(1277,-266) /sn:0 /R:14
  //: /line:"Write_Enable"
  //: /end
  //: LED g114 (w36) @(1668,-218) /sn:0 /R:3 /w:[ 3 ] /type:1
  //: joint g19 (w0) @(186, 309) /w:[ 2 -1 1 8 ]
  _GGNBUF #(2) g78 (.I(w57), .Z(w59));   //: @(-22,-464) /sn:0 /w:[ 3 0 ]
  //: joint g125 (w37) @(-142, -47) /w:[ -1 9 10 12 ]
  _GGNBUF #(2) g113 (.I(w77), .Z(w74));   //: @(1536,-372) /sn:0 /w:[ 3 0 ]
  //: SWITCH g105 (w76) @(1339,-120) /sn:0 /R:1 /w:[ 1 ] /st:0 /dn:1
  _GGBUFIF8 #(4, 6) g100 (.Z(w10), .I(w72), .E(w70));   //: @(218,52) /sn:0 /w:[ 7 0 1 ]
  //: SWITCH g93 (w66) @(775,-368) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g63 (w17) @(337,444) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: joint g43 (w77) @(1345, -372) /w:[ 2 4 -1 1 ]
  //: frame g101 @(-412,-640) /sn:0 /wi:620 /ht:299 /tx:"Memory_Read"
  //: LED g0 (w0) @(301,337) /sn:0 /R:2 /w:[ 7 ] /type:1
  //: joint g38 (w51) @(666, -162) /w:[ 2 1 -1 4 ]
  //: joint g48 (w91) @(435, 120) /w:[ 2 1 -1 4 ]
  jump_module g37 (.JEQ_enable(w20), .JNE_enable(w56), .Jump_Unconditional_Enable(w94), .status_flag(w35), .offset_enable(w80));   //: @(-752, 362) /sz:(381, 80) /R:2 /sn:0 /p:[ Ri0>0 Ri1>0 Ri2>5 Ri3>0 Lo0<0 ]
  _GGBUFIF8 #(4, 6) g95 (.Z(w51), .I(w62), .E(w68));   //: @(880,-421) /sn:0 /w:[ 0 0 1 ]
  //: SWITCH g80 (w57) @(-57,-389) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: LED g120 (w37) @(525,624) /sn:0 /R:2 /w:[ 19 ] /type:1
  //: LED g122 (w92) @(548,489) /sn:0 /w:[ 11 ] /type:0
  //: SWITCH g76 (w58) @(-133,-400) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: joint g152 (w53) @(272, -467) /w:[ 4 -1 3 10 ]
  //: LED g75 (w53) @(126,-389) /sn:0 /R:3 /w:[ 0 ] /type:1
  _GGOR6 #(14) g44 (.I0(w91), .I1(w82), .I2(w12), .I3(w47), .I4(w16), .I5(w9), .Z(w45));   //: @(809,132) /sn:0 /w:[ 3 3 3 3 3 3 0 ]
  register_file g16 (.register_input(w2), .r7_enable(w32), .r6_enable(w31), .r5_enable(w30), .r4_enable(w29), .r3_enable(w28), .r2_enable(w11), .r1_enable(w8), .r0_enable(w7), .Register_Address(w1), .Clock_Register_File(w41), .register_file_output(w86));   //: @(754, 196) /sz:(333, 258) /sn:0 /p:[ Li0>3 Li1>1 Li2>0 Li3>0 Li4>0 Li5>0 Li6>0 Li7>0 Li8>0 Li9>5 Li10>1 Ro0<9 ]
  assign w0 = w10[2:0]; //: TAP g3 @(104,309) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: joint g47 (w92) @(577, 171) /w:[ 2 -1 8 1 ]
  //: comment g143 @(-839,-142) /sn:0
  //: /line:"STATUS FLAG CLEAR CLOCK"
  //: /end
  //: joint g90 (w66) @(774, -439) /w:[ 2 4 -1 1 ]
  program_counter g26 (.offset_enable(w80), .PC_offset(w53), .PC_Clear(w14), .Program_counter_clock(w50), .PC_out(w21));   //: @(-539, -272) /sz:(357, 80) /sn:0 /p:[ Li0>3 Li1>11 Li2>1 Li3>1 Ro0<9 ]
  //: LED g109 (w51) @(725,-227) /sn:0 /R:3 /w:[ 3 ] /type:1
  //: joint g128 (w2) @(674, 216) /w:[ 2 4 1 -1 ]
  assign w3 = w10[3]; //: TAP g2 @(104,269) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:1
  _GGNBUF #(2) g91 (.I(w66), .Z(w68));   //: @(809,-439) /sn:0 /w:[ 3 0 ]
  //: joint g23 (w53) @(120, -446) /w:[ 2 -1 12 1 ]
  //: joint g141 (w22) @(-174, -162) /w:[ -1 1 2 4 ]
  //: joint g24 (w69) @(115, -7) /w:[ 2 -1 4 1 ]
  //: LED g86 (w64) @(-183,-512) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: SWITCH g39 (w50) @(-679,-188) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: LED g104 (w2) @(621,216) /sn:0 /R:1 /w:[ 0 ] /type:1
  //: joint g127 (w37) @(-197, -106) /w:[ 3 -1 4 6 ]
  //: SWITCH g110 (w78) @(1414,-154) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:1
  _GGRAM8x8 #(10, 60, 70, 10, 10, 10) g60 (.A(w53), .D(w62), .WE(w63), .OE(w66), .CS(w67));   //: @(705,-506) /w:[ 9 1 5 5 1 ]
  _GGREG #(10, 10, 20) g29 (.Q(w35), .D(w39), .EN(w43), .CLR(w84), .CK(w44));   //: @(-549,20) /sn:0 /w:[ 5 1 0 1 1 ]
  //: joint g121 (w37) @(524, 548) /w:[ 16 -1 15 18 ]
  _GGBUFIF8 #(4, 6) g82 (.Z(w53), .I(w38), .E(w59));   //: @(49,-446) /sn:0 /w:[ 13 0 1 ]
  //: joint g18 (w3) @(213, 269) /w:[ 2 -1 1 8 ]
  //: SWITCH g94 (w63) @(695,-593) /sn:0 /R:3 /w:[ 3 ] /st:1 /dn:1
  //: joint g119 (w23) @(412, 506) /w:[ -1 5 6 8 ]
  //: joint g107 (w86) @(1187, 235) /w:[ -1 6 8 5 ]
  //: joint g50 (w82) @(453, 125) /w:[ 2 4 -1 1 ]
  _GGAND3 #(8) g133 (.I0(w6), .I1(w25), .I2(w24), .Z(w26));   //: @(912,42) /sn:0 /R:1 /w:[ 0 0 0 0 ]
  //: joint g73 (w21) @(-67, -249) /w:[ 1 2 4 -1 ]
  //: joint g68 (w21) @(-134, -249) /w:[ 5 6 8 -1 ]
  //: comment g9 @(355,266) /sn:0
  //: /line:"Imm/Register"
  //: /end
  _GGBUFIF8 #(4, 6) g102 (.Z(w60), .I(w36), .E(w74));   //: @(1576,-308) /sn:0 /R:2 /w:[ 1 5 1 ]
  //: LED g71 (w80) @(-626,-331) /sn:0 /w:[ 5 ] /type:0
  //: SWITCH g59 (w15) @(355,229) /sn:0 /w:[ 0 ] /st:1 /dn:1
  ALU g22 (.adder_enable(w49), .and_enable(w91), .divider_enable(w46), .input_1_ALU(w37), .input_2_ALU(w51), .multiplier_enable(w83), .nand_enable(w12), .nor_enable(w13), .not_enable(w47), .or_enable(w9), .subtractor_enable(w16), .xor_enable(w82), .ALU_output(w48));   //: @(546, -110) /sz:(237, 226) /sn:0 /p:[ Li0>0 Li1>0 Li2>5 Li3>0 Li4>11 Li5>0 Li6>0 Li7>0 Li8>0 Li9>0 Li10>0 Li11>5 Ro0<0 ]
  //: joint g31 (w51) @(666, -122) /w:[ 6 5 8 10 ]
  _GGNBUF #(2) g87 (.I(w69), .Z(w70));   //: @(150,-7) /sn:0 /w:[ 3 0 ]
  //: SWITCH g99 (w73) @(-42,118) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  _GGADD8 #(68, 70, 62, 64) g83 (.A(w21), .B(w65), .S(w55), .CI(w61), .CO(w64));   //: @(-256,-527) /sn:0 /R:2 /w:[ 3 1 1 0 0 ]
  _GGBUFIF #(4, 6) g36 (.Z(w44), .I(w79), .E(w22));   //: @(-634,21) /sn:0 /w:[ 0 1 3 ]
  _GGOR6 #(14) g45 (.I0(w46), .I1(w49), .I2(w83), .I3(w92), .I4(w93), .I5(w13), .Z(w54));   //: @(809,168) /sn:0 /w:[ 3 3 3 5 5 3 0 ]
  _GGBUFIF8 #(4, 6) g41 (.Z(w27), .I(w37), .E(w92));   //: @(569,548) /sn:0 /w:[ 0 17 13 ]
  //: comment g69 @(-719,-255) /sn:0
  //: /line:"PC_CLEAR_CLOCK"
  //: /end
  //: joint g138 (w92) @(755, 171) /w:[ 4 6 3 -1 ]
  //: joint g42 (w37) @(485, 550) /w:[ 14 20 13 -1 ]
  //: joint g151 (w94) @(-247, 394) /w:[ 1 2 4 -1 ]
  //: LED g66 (w10) @(-1,354) /sn:0 /R:1 /w:[ 0 ] /type:1
  //: LED g146 (w20) @(-319,364) /sn:0 /w:[ 5 ] /type:0
  //: joint g28 (w24) @(962, 148) /w:[ 4 6 3 -1 ]
  //: SWITCH g34 (w40) @(-679,-132) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: joint g46 (w93) @(695, 179) /w:[ -1 2 1 8 ]
  //: joint g57 (w46) @(530, 156) /w:[ 2 4 -1 1 ]
  //: joint g150 (w56) @(-298, 410) /w:[ 2 4 1 -1 ]
  //: frame g118 @(1290,-454) /sn:0 /wi:426 /ht:372 /tx:"RAM_WRITE"
  //: DIP g84 (w65) @(-339,-458) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:1
  //: joint g14 (w0) @(301, 312) /w:[ 4 3 -1 6 ]
  _GGNBUF #(2) g11 (.I(w3), .Z(w23));   //: @(372,296) /sn:0 /w:[ 7 0 ]
  assign w4 = w10[7:4]; //: TAP g5 @(104,208) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:1
  //: LED g112 (w23) @(378,507) /sn:0 /R:1 /w:[ 7 ] /type:0
  //: joint g21 (w23) @(412, 296) /w:[ 2 -1 1 4 ]
  _GGADD8 #(68, 70, 62, 64) g61 (.A(w34), .B(w5), .S(w18), .CI(w17), .CO(w42));   //: @(309,496) /sn:0 /R:1 /w:[ 0 1 0 1 1 ]
  //: joint g123 (w92) @(576, 490) /w:[ -1 9 10 12 ]
  //: joint g32 (w37) @(-142, -107) /w:[ 1 -1 2 8 ]
  _GGMUX2x8 #(8, 8) g20 (.I0(w18), .I1(w86), .S(w23), .Z(w37));   //: @(485,519) /sn:0 /w:[ 1 0 9 21 ] /ss:0 /do:0
  //: comment g115 @(1614,-286) /sn:0 /R:14
  //: /line:"Value_to_Write"
  //: /end
  //: joint g79 (w52) @(-126, -565) /w:[ -1 1 2 4 ]
  //: joint g145 (w35) @(-549, 112) /w:[ 2 4 -1 1 ]
  //: SWITCH g97 (w71) @(129,-72) /sn:0 /R:3 /w:[ 1 ] /st:1 /dn:1
  //: joint g134 (w24) @(939, 148) /w:[ 2 1 8 -1 ]
  //: LED g148 (w94) @(-247,357) /sn:0 /w:[ 3 ] /type:0
  //: joint g129 (w1) @(500, 312) /w:[ 2 -1 1 4 ]
  //: SWITCH g89 (w67) @(697,-385) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  _GGDECODER8 #(6, 6) g15 (.I(w1), .E(w24), .Z0(w7), .Z1(w8), .Z2(w11), .Z3(w28), .Z4(w29), .Z5(w30), .Z6(w31), .Z7(w32));   //: @(546,320) /sn:0 /R:1 /w:[ 3 5 1 1 1 1 1 1 1 0 ] /ss:0 /do:0
  //: LED g147 (w56) @(-298,363) /sn:0 /w:[ 5 ] /type:0
  //: joint g27 (w53) @(342, -467) /w:[ 6 8 5 -1 ]
  //: DIP g62 (w5) @(127,483) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: frame g88 @(622,-619) /sn:0 /wi:340 /ht:270 /tx:"RAM_READ"
  //: joint g55 (w16) @(509, 140) /w:[ 2 1 -1 4 ]
  _GGMUX2x8 #(8, 8) g139 (.I0(w27), .I1(w48), .S(w26), .Z(w36));   //: @(1137,-36) /sn:0 /R:1 /w:[ 1 1 1 0 ] /ss:0 /do:0
  _GGNBUF #(2) g135 (.I(w92), .Z(w6));   //: @(849,80) /sn:0 /w:[ 7 1 ]
  _GGDECODER16 #(6, 6) g13 (.I(w4), .E(w15), .Z0(w93), .Z1(w92), .Z2(w91), .Z3(w9), .Z4(w82), .Z5(w12), .Z6(w13), .Z7(w47), .Z8(w49), .Z9(w16), .Z10(w83), .Z11(w46), .Z12(w22), .Z13(w94), .Z14(w20), .Z15(w56));   //: @(394,199) /sn:0 /R:1 /w:[ 3 1 0 0 5 5 0 5 5 5 5 5 5 0 0 0 3 3 ] /ss:0 /do:1
  //: joint g53 (w47) @(488, 143) /w:[ 2 1 -1 4 ]
  //: joint g140 (w93) @(689, 197) /w:[ 9 -1 10 12 ]

endmodule
//: /netlistEnd

//: /netlistBegin not_gate
module not_gate(not_enable, not_gate_output, not_gate_input);
//: interface  /sz:(243, 48) /bd:[ Li0>not_enable(32/48) Li1>not_gate_input[7:0](16/48) Ro0<not_gate_output[7:0](16/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [7:0] not_gate_output;    //: {0}(#:327,171)(451,171)(451,173)(50:466,173){1}
input [7:0] not_gate_input;    //: /sn:0 {0}(#:144,166)(#:169,166)(169,169)(225,169){1}
input not_enable;    //: {0}(233,164)(233,97)(234,97)(-99:234,82){1}
wire [7:0] w0;    //: /sn:0 {0}(#:241,169)(264,169)(264,171)(#:311,171){1}
//: enddecls

  //: IN g4 (not_enable) @(234,80) /sn:0 /R:3 /w:[ 1 ]
  _GGBUFIF8 #(4, 6) g3 (.Z(w0), .I(not_gate_input), .E(not_enable));   //: @(231,169) /sn:0 /w:[ 0 1 0 ]
  //: OUT g2 (not_gate_output) @(463,173) /sn:0 /w:[ 1 ]
  //: IN g1 (not_gate_input) @(142,166) /sn:0 /w:[ 0 ]
  _GGNBUF8 #(2) g0 (.I(w0), .Z(not_gate_output));   //: @(317,171) /sn:0 /w:[ 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin or_gate
module or_gate(or_gate_output, or_gate_input_2, or_gate_input_1, or_enable);
//: interface  /sz:(237, 64) /bd:[ Li0>or_enable(48/64) Li1>or_gate_input_2[7:0](32/64) Li2>or_gate_input_1[7:0](16/64) Ro0<or_gate_output[7:0](16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [7:0] or_gate_output;    //: {0}(#:357,176)(50:511,176){1}
input or_enable;    //: /sn:0 {0}(227,207)(68,207)(68,171){1}
//: {2}(68,167)(68,158)(248,158)(248,143)(238,143){3}
//: {4}(66,169)(53,169){5}
input [7:0] or_gate_input_1;    //: /sn:0 {0}(#:203,117)(233,117)(233,135){1}
input [7:0] or_gate_input_2;    //: /sn:0 {0}(232,215)(#:232,253)(#:208,253){1}
wire [7:0] w0;    //: /sn:0 {0}(#:233,151)(233,173)(336,173){1}
wire [7:0] w1;    //: /sn:0 {0}(#:232,199)(232,178)(336,178){1}
//: enddecls

  _GGBUFIF8 #(4, 6) g4 (.Z(w0), .I(or_gate_input_1), .E(or_enable));   //: @(233,141) /sn:0 /R:3 /w:[ 0 1 3 ]
  //: OUT g3 (or_gate_output) @(508,176) /sn:0 /w:[ 1 ]
  //: IN g2 (or_gate_input_2) @(206,253) /sn:0 /w:[ 1 ]
  //: IN g1 (or_gate_input_1) @(201,117) /sn:0 /w:[ 0 ]
  //: IN g6 (or_enable) @(51,169) /sn:0 /w:[ 5 ]
  //: joint g7 (or_enable) @(68, 169) /w:[ -1 2 4 1 ]
  _GGBUFIF8 #(4, 6) g5 (.Z(w1), .I(or_gate_input_2), .E(or_enable));   //: @(232,209) /sn:0 /R:1 /w:[ 0 0 0 ]
  _GGOR2x8 #(6) g0 (.I0(w0), .I1(w1), .Z(or_gate_output));   //: @(347,176) /sn:0 /w:[ 1 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin nor_gate
module nor_gate(nor_gate_output, nor_gate_input_2, nor_gate_input_1, nor_enable);
//: interface  /sz:(255, 64) /bd:[ Li0>nor_enable(48/64) Li1>nor_gate_input_2[7:0](32/64) Li2>nor_gate_input_1[7:0](16/64) Ro0<nor_gate_output[7:0](16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] nor_gate_input_2;    //: /sn:0 {0}(231,212)(#:231,250)(#:204,250){1}
output [7:0] nor_gate_output;    //: {0}(#:353,172)(374,172)(374,173)(50:507,173){1}
input [7:0] nor_gate_input_1;    //: /sn:0 {0}(231,126)(231,114)(#:199,114){1}
input nor_enable;    //: {0}(48,173)(209,173){1}
//: {2}(211,171)(211,149)(246,149)(246,134)(236,134){3}
//: {4}(211,175)(50:211,204)(226,204){5}
wire [7:0] w0;    //: /sn:0 {0}(#:231,142)(231,169)(#:50:332,169){1}
wire [7:0] w2;    //: /sn:0 {0}(#:231,196)(231,174)(#:332,174){1}
//: enddecls

  _GGBUFIF8 #(4, 6) g4 (.Z(w2), .I(nor_gate_input_2), .E(nor_enable));   //: @(231,206) /sn:0 /R:1 /w:[ 0 0 5 ]
  //: OUT g3 (nor_gate_output) @(504,173) /sn:0 /w:[ 1 ]
  //: IN g2 (nor_gate_input_2) @(202,250) /sn:0 /w:[ 1 ]
  //: IN g1 (nor_gate_input_1) @(197,114) /sn:0 /w:[ 1 ]
  //: IN g6 (nor_enable) @(46,173) /sn:0 /w:[ 0 ]
  //: joint g7 (nor_enable) @(211, 173) /w:[ -1 2 1 4 ]
  _GGBUFIF8 #(4, 6) g5 (.Z(w0), .I(nor_gate_input_1), .E(nor_enable));   //: @(231,132) /sn:0 /R:3 /w:[ 0 0 3 ]
  _GGNOR2x8 #(4) g0 (.I0(w0), .I1(w2), .Z(nor_gate_output));   //: @(343,172) /sn:0 /w:[ 1 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin ram_read
module ram_read(w6, pc_address);
//: interface  /sz:(183, 40) /bd:[ Li0>pc_address[7:0](16/40) Ro0<w6[7:0](16/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [7:0] w6;    //: /sn:0 {0}(#:758,504)(710,504)(710,486){1}
//: {2}(710,482)(#:710,477){3}
//: {4}(708,484)(698,484)(698,440)(#:684,440)(684,380)(#:606,380){5}
reg w25;    //: /sn:0 {0}(421,254)(421,259){1}
//: {2}(419,261)(409,261)(409,153){3}
//: {4}(421,263)(421,271){5}
input [7:0] pc_address;    //: /sn:0 {0}(#:184,149)(249,149)(249,296)(403,296){1}
reg w29;    //: /sn:0 {0}(346,422)(346,336)(414,336)(414,321){1}
reg w2;    //: /sn:0 {0}(490,444)(490,364){1}
//: {2}(492,362)(519,362){3}
//: {4}(490,360)(490,340)(428,340)(428,321){5}
wire [7:0] w1;    //: /sn:0 {0}(590,380)(558,380)(#:558,304)(469,304)(469,294)(#:438,294){1}
wire w28;    //: /sn:0 {0}(535,362)(598,362)(598,375){1}
//: enddecls

  //: OUT g4 (w6) @(755,504) /sn:0 /w:[ 0 ]
  _GGRAM8x8 #(10, 60, 70, 10, 10, 10) g26 (.A(pc_address), .D(w1), .WE(w25), .OE(w2), .CS(w29));   //: @(421,295) /w:[ 1 1 5 5 1 ]
  //: IN g1 (pc_address) @(182,149) /sn:0 /w:[ 0 ]
  //: SWITCH g24 (w29) @(346,436) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: joint g25 (w2) @(490, 362) /w:[ 2 4 -1 1 ]
  _GGNBUF #(2) g22 (.I(w2), .Z(w28));   //: @(525,362) /sn:0 /w:[ 3 0 ]
  //: joint g12 (w25) @(421, 261) /w:[ -1 1 2 4 ]
  //: SWITCH g11 (w2) @(490,458) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g14 (w25) @(409,140) /sn:0 /R:3 /w:[ 3 ] /st:1 /dn:1
  _GGBUFIF8 #(4, 6) g21 (.Z(w6), .I(w1), .E(w28));   //: @(596,380) /sn:0 /w:[ 5 0 1 ]
  //: joint g0 (w6) @(710, 484) /w:[ -1 2 4 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin add
module add(adder_input_2, adder_input_1, adder_enable, adder_output);
//: interface  /sz:(189, 64) /bd:[ Li0>adder_enable(48/64) Li1>adder_input_2[7:0](32/64) Li2>adder_input_1[7:0](16/64) Ro0<adder_output[7:0](16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] adder_input_1;    //: /sn:0 {0}(338,80)(338,60)(#:294,60){1}
input [7:0] adder_input_2;    //: {0}(450,75)(450,47)(#:-1:511,47){1}
reg w1;    //: /sn:0 {0}(391,203)(492,203)(492,206)(507,206){1}
input adder_enable;    //: /sn:0 {0}(343,88)(396,88)(396,83){1}
//: {2}(398,81)(408,81)(408,68)(465,68)(465,83)(455,83){3}
//: {4}(396,79)(396,25)(384,25){5}
output [7:0] adder_output;    //: {0}(#:386,327)(386,311){1}
//: {2}(388,309)(50:483,309){3}
//: {4}(386,307)(386,258)(#:367,258)(#:367,218){5}
wire w4;    //: /sn:0 {0}(218,207)(328,207)(328,203)(343,203){1}
wire [7:0] w0;    //: /sn:0 {0}(#:338,96)(338,174)(351,174)(351,189){1}
wire [7:0] w2;    //: /sn:0 {0}(#:450,91)(450,102)(460,102)(460,174)(383,174)(383,189){1}
//: enddecls

  _GGBUFIF8 #(4, 6) g8 (.Z(w0), .I(adder_input_1), .E(adder_enable));   //: @(338,86) /sn:0 /R:3 /w:[ 0 0 0 ]
  //: SWITCH g4 (w1) @(525,206) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  //: LED g3 (adder_output) @(386,334) /sn:0 /R:2 /w:[ 0 ] /type:1
  //: IN g2 (adder_input_2) @(513,47) /sn:0 /R:2 /w:[ 1 ]
  //: IN g1 (adder_input_1) @(292,60) /sn:0 /w:[ 1 ]
  //: IN g10 (adder_enable) @(382,25) /sn:0 /w:[ 5 ]
  //: OUT g6 (adder_output) @(480,309) /sn:0 /w:[ 3 ]
  _GGBUFIF8 #(4, 6) g9 (.Z(w2), .I(adder_input_2), .E(adder_enable));   //: @(450,81) /sn:0 /R:3 /w:[ 0 0 3 ]
  //: joint g7 (adder_output) @(386, 309) /w:[ 2 4 -1 1 ]
  //: joint g11 (adder_enable) @(396, 81) /w:[ 2 4 -1 1 ]
  //: LED g5 (w4) @(211,207) /sn:0 /R:1 /w:[ 0 ] /type:0
  _GGADD8 #(68, 70, 62, 64) g0 (.A(w0), .B(w2), .S(adder_output), .CI(w1), .CO(w4));   //: @(367,205) /sn:0 /w:[ 1 1 5 0 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin and_gate
module and_gate(and_gate_output, and_gate_input_2, and_gate_input_1, and_enable);
//: interface  /sz:(255, 64) /bd:[ Li0>and_enable(48/64) Li1>and_gate_input_2[7:0](32/64) Li2>and_gate_input_1[7:0](16/64) Ro0<and_gate_output[7:0](16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [7:0] and_gate_output;    //: {0}(#:368,188)(50:516,188){1}
input [7:0] and_gate_input_1;    //: /sn:0 {0}(229,136)(229,129)(#:208,129){1}
input and_enable;    //: {0}(60,190)(206,190){1}
//: {2}(208,188)(208,159)(244,159)(244,144)(234,144){3}
//: {4}(208,192)(50:208,224)(223,224){5}
input [7:0] and_gate_input_2;    //: /sn:0 {0}(228,232)(#:228,265)(#:213,265){1}
wire [7:0] w0;    //: /sn:0 {0}(#:229,152)(229,185)(#:347,185){1}
wire [7:0] w1;    //: /sn:0 {0}(#:228,216)(228,190)(#:347,190){1}
//: enddecls

  _GGBUFIF8 #(4, 6) g4 (.Z(w0), .I(and_gate_input_1), .E(and_enable));   //: @(229,142) /sn:0 /R:3 /w:[ 0 0 3 ]
  //: OUT g3 (and_gate_output) @(513,188) /sn:0 /w:[ 1 ]
  //: IN g2 (and_gate_input_2) @(211,265) /sn:0 /w:[ 1 ]
  //: IN g1 (and_gate_input_1) @(206,129) /sn:0 /w:[ 1 ]
  //: IN g6 (and_enable) @(58,190) /sn:0 /w:[ 0 ]
  //: joint g7 (and_enable) @(208, 190) /w:[ -1 2 1 4 ]
  _GGBUFIF8 #(4, 6) g5 (.Z(w1), .I(and_gate_input_2), .E(and_enable));   //: @(228,226) /sn:0 /R:1 /w:[ 0 0 5 ]
  _GGAND2x8 #(6) g0 (.I0(w0), .I1(w1), .Z(and_gate_output));   //: @(358,188) /sn:0 /w:[ 1 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin subtractor
module subtractor(subtractor_out, to_be_subtracted, subtractor_input_2, subtractor_enable);
//: interface  /sz:(291, 64) /bd:[ Li0>subtractor_enable(48/64) Li1>to_be_subtracted[7:0](32/64) Li2>subtractor_input_2[7:0](16/64) Ro0<subtractor_out[7:0](16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [7:0] subtractor_out;    //: {0}(#:50:493,344)(387,344){1}
//: {2}(385,342)(#:385,266){3}
//: {4}(#:383,344)(301,344)(301,329){5}
input subtractor_enable;    //: /sn:0 {0}(315,140)(369,140){1}
//: {2}(371,138)(371,33){3}
//: {4}(371,142)(371,145)(416,145)(416,160)(406,160){5}
input [7:0] to_be_subtracted;    //: /sn:0 {0}(310,132)(310,125)(#:245,125){1}
reg w1;    //: /sn:0 {0}(409,251)(489,251)(489,248)(504,248){1}
input [7:0] subtractor_input_2;    //: {0}(401,152)(401,133)(#:-99:488,133){1}
wire w4;    //: /sn:0 {0}(276,259)(346,259)(346,251)(361,251){1}
wire [7:0] w3;    //: /sn:0 {0}(#:401,168)(401,237){1}
wire [7:0] w0;    //: /sn:0 {0}(#:344,182)(369,182)(369,237){1}
wire [7:0] w2;    //: /sn:0 {0}(#:310,148)(310,182)(328,182){1}
//: enddecls

  //: joint g8 (subtractor_out) @(385, 344) /w:[ 1 2 4 -1 ]
  //: OUT g4 (subtractor_out) @(490,344) /sn:0 /w:[ 0 ]
  //: IN g3 (to_be_subtracted) @(243,125) /sn:0 /w:[ 1 ]
  //: IN g2 (subtractor_input_2) @(490,133) /sn:0 /R:2 /w:[ 1 ]
  _GGNBUF8 #(2) g1 (.I(w2), .Z(w0));   //: @(334,182) /sn:0 /w:[ 1 0 ]
  _GGBUFIF8 #(4, 6) g10 (.Z(w3), .I(subtractor_input_2), .E(subtractor_enable));   //: @(401,158) /sn:0 /R:3 /w:[ 0 0 5 ]
  //: LED g6 (w4) @(269,259) /sn:0 /R:1 /w:[ 0 ] /type:0
  _GGBUFIF8 #(4, 6) g9 (.Z(w2), .I(to_be_subtracted), .E(subtractor_enable));   //: @(310,138) /sn:0 /R:3 /w:[ 0 0 0 ]
  //: LED g7 (subtractor_out) @(301,322) /sn:0 /w:[ 5 ] /type:1
  //: joint g12 (subtractor_enable) @(371, 140) /w:[ -1 2 1 4 ]
  //: IN g11 (subtractor_enable) @(371,31) /sn:0 /R:3 /w:[ 3 ]
  //: SWITCH g5 (w1) @(522,248) /sn:0 /R:2 /w:[ 1 ] /st:1 /dn:1
  _GGADD8 #(68, 70, 62, 64) g0 (.A(w0), .B(w3), .S(subtractor_out), .CI(w1), .CO(w4));   //: @(385,253) /sn:0 /w:[ 1 1 3 0 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin divider
module divider(divider_output, divider_input_2, divider_input_register, divider_enable);
//: interface  /sz:(321, 64) /bd:[ Li0>divider_enable(48/64) Li1>divider_input_register[7:0](32/64) Li2>divider_input_2[7:0](16/64) Ro0<divider_output[7:0](16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input divider_enable;    //: {0}(327,68)(327,43)(354,43){1}
//: {2}(358,43)(410,43)(410,86)(423,86)(423,76){3}
//: {4}(356,41)(-86:356,28){5}
input [7:0] divider_input_2;    //: /sn:0 {0}(431,71)(475,71)(#:475,72)(#:542,72){1}
output [7:0] divider_output;    //: {0}(#:367,186)(367,239)(379,239){1}
//: {2}(383,239)(50:480,239){3}
//: {4}(381,241)(#:381,251)(382,251)(382,265){5}
input [7:0] divider_input_register;    //: /sn:0 {0}(#:264,76)(304,76)(304,73)(319,73){1}
wire [7:0] w0;    //: /sn:0 {0}(#:415,71)(373,71)(#:373,157){1}
wire [7:0] w3;    //: /sn:0 {0}(230,240)(347,240)(#:347,186){1}
wire [7:0] w1;    //: /sn:0 {0}(#:335,73)(341,73)(#:341,157){1}
//: enddecls

  _GGBUFIF8 #(4, 6) g8 (.Z(w0), .I(divider_input_2), .E(divider_enable));   //: @(425,71) /sn:0 /R:2 /w:[ 0 0 3 ]
  //: OUT g4 (divider_output) @(477,239) /sn:0 /w:[ 3 ]
  //: LED g3 (w3) @(223,240) /sn:0 /R:1 /w:[ 0 ] /type:1
  //: IN g2 (divider_input_2) @(544,72) /sn:0 /R:2 /w:[ 1 ]
  //: IN g1 (divider_input_register) @(262,76) /sn:0 /w:[ 0 ]
  //: joint g10 (divider_enable) @(356, 43) /w:[ 2 4 1 -1 ]
  //: joint g6 (divider_output) @(381, 239) /w:[ 2 -1 1 4 ]
  //: IN g9 (divider_enable) @(356,26) /sn:0 /R:3 /w:[ 5 ]
  _GGBUFIF8 #(4, 6) g7 (.Z(w1), .I(divider_input_register), .E(divider_enable));   //: @(325,73) /sn:0 /w:[ 0 1 0 ]
  //: LED g5 (divider_output) @(382,272) /sn:0 /R:2 /w:[ 5 ] /type:1
  _GGDIV8 #(236, 236) g0 (.A(w1), .B(w0), .Q(divider_output), .R(w3));   //: @(357,173) /sn:0 /w:[ 1 1 0 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin nand_gate
module nand_gate(nand_gate_output, nand_gate_input_2, nand_gate_input_1, nand_enable);
//: interface  /sz:(273, 64) /bd:[ Li0>nand_enable(48/64) Li1>nand_gate_input_2[7:0](32/64) Li2>nand_gate_input_1[7:0](16/64) Ro0<nand_gate_output[7:0](16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] nand_gate_input_2;    //: /sn:0 {0}(236,215)(236,237)(#:226,237)(#:226,255)(#:211,255){1}
input [7:0] nand_gate_input_1;    //: /sn:0 {0}(234,133)(#:234,98)(225,98)(225,119)(#:206,119){1}
input nand_enable;    //: /sn:0 {0}(231,207)(162,207)(162,190){1}
//: {2}(162,186)(162,156)(249,156)(249,141)(239,141){3}
//: {4}(160,188)(147,188){5}
output [7:0] nand_gate_output;    //: {0}(#:353,177)(378,177)(99:378,178)(514,178){1}
wire [7:0] w0;    //: /sn:0 {0}(#:50:332,174)(234,174)(#:234,149){1}
wire [7:0] w1;    //: /sn:0 {0}(#:236,199)(236,179)(#:50:332,179){1}
//: enddecls

  _GGBUFIF8 #(4, 6) g4 (.Z(w0), .I(nand_gate_input_1), .E(nand_enable));   //: @(234,139) /sn:0 /R:3 /w:[ 1 0 3 ]
  //: OUT g3 (nand_gate_output) @(511,178) /sn:0 /w:[ 1 ]
  //: IN g2 (nand_gate_input_2) @(209,255) /sn:0 /w:[ 1 ]
  //: IN g1 (nand_gate_input_1) @(204,119) /sn:0 /w:[ 1 ]
  //: IN g6 (nand_enable) @(145,188) /sn:0 /w:[ 5 ]
  //: joint g7 (nand_enable) @(162, 188) /w:[ -1 2 4 1 ]
  _GGBUFIF8 #(4, 6) g5 (.Z(w1), .I(nand_gate_input_2), .E(nand_enable));   //: @(236,209) /sn:0 /R:1 /w:[ 0 0 0 ]
  _GGNAND2x8 #(4) g0 (.I0(w0), .I1(w1), .Z(nand_gate_output));   //: @(343,177) /sn:0 /w:[ 0 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU
module ALU(adder_enable, subtractor_enable, input_2_ALU, multiplier_enable, and_enable, xor_enable, nand_enable, or_enable, divider_enable, input_1_ALU, ALU_output, not_enable, nor_enable);
//: interface  /sz:(237, 230) /bd:[ Li0>input_1_ALU[7:0](3/230) Li1>input_2_ALU[7:0](14/230) Li2>and_enable(25/230) Li3>or_enable(37/230) Li4>xor_enable(49/230) Li5>nand_enable(67/230) Li6>nor_enable(85/230) Li7>not_enable(109/230) Li8>adder_enable(135/230) Li9>subtractor_enable(157/230) Li10>multiplier_enable(173/230) Li11>divider_enable(214/230) Ro0<ALU_output[7:0](17/230) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input multiplier_enable;    //: /sn:0 {0}(163,238)(141,238){1}
//: {2}(139,236)(139,235)(81,235){3}
//: {4}(137,238)(127,238)(127,223)(492,223)(492,192)(507,192)(507,202){5}
input divider_enable;    //: {0}(163,380)(145,380)(145,425){1}
//: {2}(147,427)(527,427)(527,336)(537,336)(537,346){3}
//: {4}(145,429)(-99:145,461){5}
input [7:0] input_1_ALU;    //: /sn:0 {0}(#:163,-68)(114,-68)(114,-74){1}
//: {2}(116,-76)(#:126,-76)(126,68){3}
//: {4}(128,70)(163,70){5}
//: {6}(#:126,72)(126,193){7}
//: {8}(128,195)(#:138,195)(138,364)(163,364){9}
//: {10}(126,197)(126,206)(163,206){11}
//: {12}(114,-78)(#:114,-129)(-325,-129){13}
//: {14}(-327,-131)(#:-327,-168){15}
//: {16}(#:-327,-127)(-327,-88){17}
//: {18}(-325,-86)(-271,-86)(-271,-87)(-217,-87){19}
//: {20}(#:-327,-84)(-327,19){21}
//: {22}(-325,21)(#:-315,21)(-315,150){23}
//: {24}(-313,152)(-217,152){25}
//: {26}(#:-315,154)(-315,298){27}
//: {28}(-313,300)(-222,300){29}
//: {30}(#:-315,302)(-315,395)(-224,395){31}
//: {32}(-327,23)(-327,25)(-217,25){33}
input xor_enable;    //: {0}(-353,181)(-284,181){1}
//: {2}(-280,181)(-230,181)(50:-230,184)(-217,184){3}
//: {4}(-282,179)(-282,169)(72,169)(72,180){5}
output [7:0] ALU_output;    //: {0}(#:82,513)(659,513)(659,423){1}
//: {2}(659,419)(659,358){3}
//: {4}(659,354)(659,325){5}
//: {6}(659,321)(659,245){7}
//: {8}(661,243)(#:671,243)(671,242)(50:821,242){9}
//: {10}(659,241)(659,212){11}
//: {12}(659,208)(659,185){13}
//: {14}(659,181)(659,49){15}
//: {16}(659,45)(659,23){17}
//: {18}(659,19)(659,-34){19}
//: {20}(659,-38)(659,-68)(#:409,-68){21}
//: {22}(657,-36)(#:78,-36){23}
//: {24}(657,21)(648,21)(648,10)(#:66,10){25}
//: {26}(657,47)(647,47)(647,51)(#:510,51){27}
//: {28}(657,183)(647,183)(647,185)(#:80,185){29}
//: {30}(657,210)(647,210)(647,207)(#:515,207){31}
//: {32}(657,323)(647,323)(647,325)(#:73,325){33}
//: {34}(657,356)(647,356)(647,351)(#:545,351){35}
//: {36}(657,421)(#:93,421){37}
input or_enable;    //: /sn:0 {0}(-217,57)(-240,57){1}
//: {2}(-242,55)(-242,-2)(58,-2)(58,5){3}
//: {4}(-244,57)(-314,57)(-314,58)(-327,58){5}
input subtractor_enable;    //: {0}(163,86)(154,86)(-97:154,88)(137,88){1}
//: {2}(135,86)(135,76)(487,76)(487,36)(502,36)(502,46){3}
//: {4}(133,88)(77,88){5}
input and_enable;    //: /sn:0 {0}(-217,-55)(-272,-55){1}
//: {2}(-276,-55)(-319,-55)(-319,-53)(-332,-53){3}
//: {4}(-274,-53)(-274,-51)(70,-51)(70,-41){5}
input adder_enable;    //: /sn:0 {0}(163,-36)(130,-36)(130,-138){1}
//: {2}(132,-140)(401,-140)(401,-73){3}
//: {4}(130,-142)(130,-161){5}
input not_enable;    //: /sn:0 {0}(-217,526)(-280,526){1}
//: {2}(-282,524)(-282,514)(59,514)(59,498)(74,498)(74,508){3}
//: {4}(-284,526)(-360,526){5}
input [7:0] input_2_ALU;    //: {0}(#:-99:-417,571)(-298,571){1}
//: {2}(-294,571)(-239,571){3}
//: {4}(-235,571)(152,571){5}
//: {6}(156,571)(191,571)(191,559){7}
//: {8}(#:154,569)(154,410)(109,410)(109,350){9}
//: {10}(111,348)(163,348){11}
//: {12}(#:109,346)(109,224){13}
//: {14}(111,222)(163,222){15}
//: {16}(#:109,220)(109,118)(109,118)(109,56){17}
//: {18}(111,54)(163,54){19}
//: {20}(#:109,52)(109,-52)(163,-52){21}
//: {22}(#:-237,569)(-237,512){23}
//: {24}(-235,510)(-217,510){25}
//: {26}(#:-237,508)(-237,418){27}
//: {28}(-237,414)(-237,411)(-224,411){29}
//: {30}(-239,416)(#:-265,416)(-265,316)(-242,316){31}
//: {32}(-238,316)(-222,316){33}
//: {34}(#:-240,314)(-240,176){35}
//: {36}(-240,172)(-240,168)(-217,168){37}
//: {38}(-242,174)(#:-261,174)(-261,41)(-217,41){39}
//: {40}(#:-296,569)(-296,-71)(-217,-71){41}
input nor_enable;    //: /sn:0 {0}(-222,332)(-247,332){1}
//: {2}(-249,330)(-249,310)(65,310)(65,320){3}
//: {4}(-251,332)(-337,332)(-337,316)(-345,316){5}
input nand_enable;    //: {0}(-349,425)(-270,425){1}
//: {2}(-266,425)(-237,425)(50:-237,427)(-224,427){3}
//: {4}(-268,423)(-268,413)(85,413)(85,416){5}
wire [7:0] w7;    //: /sn:0 {0}(529,351)(504,351)(#:504,348)(486,348){1}
wire [7:0] w34;    //: /sn:0 {0}(494,51)(471,51)(#:471,54)(456,54){1}
wire [7:0] w0;    //: /sn:0 {0}(#:393,-68)(354,-68){1}
wire [7:0] w3;    //: /sn:0 {0}(#:67,-87)(53,-87){1}
//: {2}(49,-87)(40,-87){3}
//: {4}(#:51,-85)(51,-36)(62,-36){5}
wire [7:0] w30;    //: /sn:0 {0}(66,513)(38,513)(#:38,510)(28,510){1}
wire [7:0] w19;    //: /sn:0 {0}(#:65,152)(51,152){1}
//: {2}(47,152)(40,152){3}
//: {4}(#:49,154)(49,185)(64,185){5}
wire [7:0] w23;    //: /sn:0 {0}(#:51,300)(44,300){1}
//: {2}(40,300)(35,300){3}
//: {4}(#:42,302)(42,325)(57,325){5}
wire [7:0] w27;    //: /sn:0 {0}(77,421)(62,421)(#:62,395)(51,395){1}
wire [7:0] w15;    //: /sn:0 {0}(#:58,25)(37,25){1}
//: {2}(#:35,23)(35,10)(50,10){3}
//: {4}(33,25)(22,25){5}
wire [7:0] w38;    //: /sn:0 {0}(499,207)(479,207)(#:479,206)(468,206){1}
//: enddecls

  subtractor g8 (.subtractor_input_2(input_2_ALU), .to_be_subtracted(input_1_ALU), .subtractor_enable(subtractor_enable), .subtractor_out(w34));   //: @(164, 38) /sz:(291, 64) /sn:0 /p:[ Li0>19 Li1>5 Li2>0 Ro0<1 ]
  xor_gate g4 (.xor_gate_input_1(input_1_ALU), .xor_gate_input_2(input_2_ALU), .xor_enable(xor_enable), .xor_gate_output(w19));   //: @(-216, 136) /sz:(255, 64) /sn:0 /p:[ Li0>25 Li1>37 Li2>3 Ro0<3 ]
  _GGBUFIF8 #(4, 6) g44 (.Z(ALU_output), .I(w34), .E(subtractor_enable));   //: @(500,51) /sn:0 /w:[ 27 0 3 ]
  //: IN g16 (adder_enable) @(130,-163) /sn:0 /R:3 /w:[ 5 ]
  or_gate g3 (.or_gate_input_1(input_1_ALU), .or_gate_input_2(input_2_ALU), .or_enable(or_enable), .or_gate_output(w15));   //: @(-216, 9) /sz:(237, 64) /sn:0 /p:[ Li0>33 Li1>39 Li2>0 Ro0<5 ]
  //: joint g47 (multiplier_enable) @(139, 238) /w:[ 1 2 4 -1 ]
  //: joint g26 (input_1_ALU) @(114, -76) /w:[ 2 12 -1 1 ]
  //: IN g17 (subtractor_enable) @(75,88) /sn:0 /w:[ 5 ]
  and_gate g2 (.and_gate_input_1(input_1_ALU), .and_gate_input_2(input_2_ALU), .and_enable(and_enable), .and_gate_output(w3));   //: @(-216, -103) /sz:(255, 64) /sn:0 /p:[ Li0>19 Li1>41 Li2>0 Ro0<3 ]
  //: joint g30 (input_2_ALU) @(-296, 571) /w:[ 2 40 1 -1 ]
  //: joint g23 (input_1_ALU) @(-327, 21) /w:[ 22 21 -1 32 ]
  //: joint g39 (input_2_ALU) @(109, 54) /w:[ 18 20 -1 17 ]
  //: joint g24 (input_1_ALU) @(-315, 152) /w:[ 24 23 -1 26 ]
  divider g1 (.divider_input_2(input_2_ALU), .divider_input_register(input_1_ALU), .divider_enable(divider_enable), .divider_output(w7));   //: @(164, 332) /sz:(321, 64) /sn:0 /p:[ Li0>11 Li1>9 Li2>0 Ro0<1 ]
  //: IN g29 (input_2_ALU) @(-419,571) /sn:0 /w:[ 0 ]
  _GGBUFIF8 #(4, 6) g60 (.Z(ALU_output), .I(w15), .E(or_enable));   //: @(56,10) /sn:0 /w:[ 25 3 3 ]
  //: joint g51 (not_enable) @(-282, 526) /w:[ 1 2 4 -1 ]
  //: IN g18 (multiplier_enable) @(79,235) /sn:0 /w:[ 3 ]
  //: joint g70 (ALU_output) @(659, 210) /w:[ -1 12 30 11 ]
  //: joint g25 (input_1_ALU) @(-315, 300) /w:[ 28 27 -1 30 ]
  //: IN g10 (and_enable) @(-334,-53) /sn:0 /w:[ 3 ]
  //: joint g65 (and_enable) @(-274, -55) /w:[ 1 -1 2 4 ]
  //: joint g64 (w3) @(51, -87) /w:[ 1 -1 2 4 ]
  //: joint g49 (divider_enable) @(145, 427) /w:[ 2 1 -1 4 ]
  //: joint g72 (ALU_output) @(659, 323) /w:[ -1 6 32 5 ]
  nand_gate g6 (.nand_gate_input_1(input_1_ALU), .nand_gate_input_2(input_2_ALU), .nand_enable(nand_enable), .nand_gate_output(w27));   //: @(-223, 379) /sz:(273, 64) /sn:0 /p:[ Li0>31 Li1>29 Li2>3 Ro0<1 ]
  _GGBUFIF8 #(4, 6) g50 (.Z(ALU_output), .I(w30), .E(not_enable));   //: @(72,513) /sn:0 /w:[ 0 0 3 ]
  //: joint g35 (input_2_ALU) @(-240, 174) /w:[ -1 36 38 35 ]
  multiplier g9 (.multiplier_input_1(input_1_ALU), .multiplier_input_2(input_2_ALU), .multiplier_enable(multiplier_enable), .multiplier_output_1(w38));   //: @(164, 190) /sz:(303, 64) /sn:0 /p:[ Li0>11 Li1>15 Li2>0 Ro0<1 ]
  not_gate g7 (.not_gate_input(input_2_ALU), .not_enable(not_enable), .not_gate_output(w30));   //: @(-216, 494) /sz:(243, 48) /sn:0 /p:[ Li0>25 Li1>0 Ro0<1 ]
  //: joint g56 (nor_enable) @(-249, 332) /w:[ 1 2 4 -1 ]
  //: joint g58 (w19) @(49, 152) /w:[ 1 -1 2 4 ]
  //: joint g68 (ALU_output) @(659, 21) /w:[ -1 18 24 17 ]
  //: joint g73 (ALU_output) @(659, 421) /w:[ -1 2 36 1 ]
  //: joint g31 (input_2_ALU) @(-237, 571) /w:[ 4 22 3 -1 ]
  //: joint g22 (input_1_ALU) @(-327, -86) /w:[ 18 17 -1 20 ]
  //: joint g59 (xor_enable) @(-282, 181) /w:[ 2 4 1 -1 ]
  //: joint g71 (ALU_output) @(659, 356) /w:[ -1 4 34 3 ]
  //: joint g67 (ALU_output) @(659, 47) /w:[ -1 16 26 15 ]
  //: joint g36 (input_2_ALU) @(154, 571) /w:[ 6 8 5 -1 ]
  //: joint g33 (input_2_ALU) @(-237, 416) /w:[ -1 28 30 27 ]
  //: joint g41 (adder_enable) @(130, -140) /w:[ 2 4 -1 1 ]
  //: joint g45 (subtractor_enable) @(135, 88) /w:[ 1 2 4 -1 ]
  _GGBUFIF8 #(4, 6) g54 (.Z(ALU_output), .I(w23), .E(nor_enable));   //: @(63,325) /sn:0 /w:[ 33 5 3 ]
  _GGBUFIF8 #(4, 6) g40 (.Z(ALU_output), .I(w0), .E(adder_enable));   //: @(399,-68) /sn:0 /w:[ 21 0 3 ]
  _GGBUFIF8 #(4, 6) g52 (.Z(ALU_output), .I(w27), .E(nand_enable));   //: @(83,421) /sn:0 /w:[ 37 0 5 ]
  //: joint g69 (ALU_output) @(659, 183) /w:[ -1 14 28 13 ]
  //: joint g42 (ALU_output) @(659, 243) /w:[ 8 10 -1 7 ]
  //: joint g66 (ALU_output) @(659, -36) /w:[ -1 20 22 19 ]
  //: IN g12 (xor_enable) @(-355,181) /sn:0 /w:[ 0 ]
  //: joint g34 (input_2_ALU) @(-240, 316) /w:[ 32 34 31 -1 ]
  //: joint g28 (input_1_ALU) @(126, 195) /w:[ 8 7 -1 10 ]
  _GGBUFIF8 #(4, 6) g46 (.Z(ALU_output), .I(w38), .E(multiplier_enable));   //: @(505,207) /sn:0 /w:[ 31 0 5 ]
  _GGBUFIF8 #(4, 6) g57 (.Z(ALU_output), .I(w19), .E(xor_enable));   //: @(70,185) /sn:0 /w:[ 29 5 5 ]
  //: IN g14 (nand_enable) @(-351,425) /sn:0 /w:[ 0 ]
  //: IN g11 (or_enable) @(-329,58) /sn:0 /w:[ 5 ]
  nor_gate g5 (.nor_gate_input_1(input_1_ALU), .nor_gate_input_2(input_2_ALU), .nor_enable(nor_enable), .nor_gate_output(w23));   //: @(-221, 284) /sz:(255, 64) /sn:0 /p:[ Li0>29 Li1>33 Li2>0 Ro0<3 ]
  //: joint g21 (input_1_ALU) @(-327, -129) /w:[ 13 14 -1 16 ]
  //: IN g19 (divider_enable) @(145,463) /sn:0 /R:1 /w:[ 5 ]
  //: joint g61 (w15) @(35, 25) /w:[ 1 2 4 -1 ]
  //: joint g32 (input_2_ALU) @(-237, 510) /w:[ 24 26 -1 23 ]
  //: IN g20 (input_1_ALU) @(-327,-170) /sn:0 /R:3 /w:[ 15 ]
  _GGBUFIF8 #(4, 6) g63 (.Z(ALU_output), .I(w3), .E(and_enable));   //: @(68,-36) /sn:0 /w:[ 23 5 5 ]
  //: OUT g43 (ALU_output) @(818,242) /sn:0 /w:[ 9 ]
  //: joint g38 (input_2_ALU) @(109, 222) /w:[ 14 16 -1 13 ]
  //: IN g15 (not_enable) @(-362,526) /sn:0 /w:[ 5 ]
  add g0 (.adder_input_1(input_1_ALU), .adder_input_2(input_2_ALU), .adder_enable(adder_enable), .adder_output(w0));   //: @(164, -84) /sz:(189, 64) /sn:0 /p:[ Li0>0 Li1>21 Li2>0 Ro0<1 ]
  //: joint g27 (input_1_ALU) @(126, 70) /w:[ 4 3 -1 6 ]
  _GGBUFIF8 #(4, 6) g48 (.Z(ALU_output), .I(w7), .E(divider_enable));   //: @(535,351) /sn:0 /w:[ 35 0 3 ]
  //: joint g37 (input_2_ALU) @(109, 348) /w:[ 10 12 -1 9 ]
  //: joint g62 (or_enable) @(-242, 57) /w:[ 1 2 4 -1 ]
  //: joint g55 (w23) @(42, 300) /w:[ 1 -1 2 4 ]
  //: IN g13 (nor_enable) @(-347,316) /sn:0 /w:[ 5 ]
  //: joint g53 (nand_enable) @(-268, 425) /w:[ 2 4 1 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin multiplier
module multiplier(multiplier_enable, multiplier_output_1, multiplier_input_2, multiplier_input_1);
//: interface  /sz:(303, 64) /bd:[ Li0>multiplier_enable(48/64) Li1>multiplier_input_2[7:0](32/64) Li2>multiplier_input_1[7:0](16/64) Ro0<multiplier_output_1[7:0](16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input multiplier_enable;    //: /sn:0 {0}(297,85)(297,44)(349,44){1}
//: {2}(353,44)(382,44)(382,110)(395,110)(395,103){3}
//: {4}(351,42)(351,29){5}
input [7:0] multiplier_input_1;    //: /sn:0 {0}(289,90)(251,90)(#:251,83)(#:216,83){1}
input [7:0] multiplier_input_2;    //: {0}(403,98)(458,98)(#:458,106)(#:99:488,106){1}
output [7:0] multiplier_output_1;    //: {0}(#:345,200)(345,310){1}
//: {2}(347,312)(50:455,312){3}
//: {4}(#:343,312)(193,312)(193,284){5}
wire [7:0] w1;    //: /sn:0 {0}(#:305,90)(329,90)(#:329,171){1}
wire [7:0] w2;    //: /sn:0 {0}(#:387,98)(361,98)(#:361,171){1}
//: enddecls

  //: IN g8 (multiplier_enable) @(351,27) /sn:0 /R:3 /w:[ 5 ]
  //: LED g4 (multiplier_output_1) @(193,277) /sn:0 /w:[ 5 ] /type:1
  //: OUT g3 (multiplier_output_1) @(452,312) /sn:0 /w:[ 3 ]
  //: IN g2 (multiplier_input_2) @(490,106) /sn:0 /R:2 /w:[ 1 ]
  //: IN g1 (multiplier_input_1) @(214,83) /sn:0 /w:[ 1 ]
  _GGBUFIF8 #(4, 6) g6 (.Z(w1), .I(multiplier_input_1), .E(multiplier_enable));   //: @(295,90) /sn:0 /w:[ 0 0 0 ]
  //: joint g9 (multiplier_enable) @(351, 44) /w:[ 2 4 1 -1 ]
  _GGBUFIF8 #(4, 6) g7 (.Z(w2), .I(multiplier_input_2), .E(multiplier_enable));   //: @(397,98) /sn:0 /R:2 /w:[ 0 0 3 ]
  //: joint g5 (multiplier_output_1) @(345, 312) /w:[ 2 1 4 -1 ]
  _GGMUL8 #(124) g0 (.A(w1), .B(w2), .P(multiplier_output_1));   //: @(345,187) /sn:0 /w:[ 1 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin jump_module
module jump_module(JEQ_enable, JNE_enable, Jump_Unconditional_Enable, offset_enable, status_flag);
//: interface  /sz:(381, 80) /bd:[ Li0>status_flag(64/80) Li1>Jump_Unconditional_Enable(48/80) Li2>JNE_enable(32/80) Li3>JEQ_enable(16/80) Ro0<offset_enable(16/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input JNE_enable;    //: {0}(469,194)(554,194)(46:554,199)(569,199){1}
output offset_enable;    //: {0}(50:855,235)(844,235)(844,231)(715,231){1}
input Jump_Unconditional_Enable;    //: /sn:0 {0}(621,330)(688,330)(688,236)(694,236){1}
input JEQ_enable;    //: /sn:0 {0}(566,296)(441,296)(441,307)(426,307){1}
input status_flag;    //: /sn:0 {0}(569,204)(481,204)(481,243){1}
//: {2}(479,245)(466,245){3}
//: {4}(481,247)(481,277)(495,277){5}
wire w3;    //: /sn:0 {0}(511,277)(551,277)(551,291)(566,291){1}
wire w2;    //: /sn:0 {0}(590,202)(679,202)(679,226)(694,226){1}
wire w5;    //: /sn:0 {0}(587,294)(679,294)(679,231)(694,231){1}
//: enddecls

  //: IN g8 (JEQ_enable) @(424,307) /sn:0 /w:[ 1 ]
  //: IN g4 (JNE_enable) @(467,194) /sn:0 /w:[ 0 ]
  //: IN g3 (Jump_Unconditional_Enable) @(619,330) /sn:0 /w:[ 0 ]
  _GGOR3 #(8) g2 (.I0(w2), .I1(w5), .I2(Jump_Unconditional_Enable), .Z(offset_enable));   //: @(705,231) /sn:0 /w:[ 1 1 1 1 ]
  _GGAND2 #(6) g1 (.I0(w3), .I1(JEQ_enable), .Z(w5));   //: @(577,294) /sn:0 /w:[ 1 0 0 ]
  _GGNBUF #(2) g6 (.I(status_flag), .Z(w3));   //: @(501,277) /sn:0 /w:[ 5 0 ]
  //: OUT g9 (offset_enable) @(852,235) /sn:0 /w:[ 0 ]
  //: joint g7 (status_flag) @(481, 245) /w:[ -1 1 2 4 ]
  //: IN g5 (status_flag) @(464,245) /sn:0 /w:[ 3 ]
  _GGAND2 #(6) g0 (.I0(JNE_enable), .I1(status_flag), .Z(w2));   //: @(580,202) /sn:0 /w:[ 1 0 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin register_file
module register_file(register_file_output, Clock_Register_File, r7_enable, r1_enable, r0_enable, r6_enable, r2_enable, Register_Address, register_input, r5_enable, r3_enable, r4_enable);
//: interface  /sz:(333, 258) /bd:[ Li0>Clock_Register_File(242/258) Li1>Register_Address[2:0](226/258) Li2>r0_enable(206/258) Li3>r1_enable(189/258) Li4>r2_enable(169/258) Li5>r3_enable(142/258) Li6>r4_enable(115/258) Li7>r5_enable(86/258) Li8>r6_enable(64/258) Li9>r7_enable(44/258) Li10>register_input[7:0](15/258) Ro0<register_file_output[7:0](16/258) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input r5_enable;    //: /sn:0 {0}(847,342)(862,342)(862,341)(888,341){1}
output [7:0] register_file_output;    //: {0}(#:1172,356)(1210,356)(1210,417)(1203,417)(1203,432)(50:1213,432){1}
input r4_enable;    //: /sn:0 {0}(849,418)(888,418)(888,419)(901,419){1}
input r2_enable;    //: /sn:0 {0}(854,553)(880,553){1}
input r1_enable;    //: /sn:0 {0}(848,623)(878,623)(878,626)(890,626){1}
input [7:0] register_input;    //: {0}(#:597,92)(612,92){1}
//: {2}(#:616,92)(714,92)(714,182){3}
//: {4}(99:614,94)(614,242){5}
//: {6}(#:616,244)(714,244)(714,258){7}
//: {8}(614,246)(614,301){9}
//: {10}(#:616,303)(714,303)(714,326){11}
//: {12}(614,305)(614,375){13}
//: {14}(#:616,377)(714,377)(714,393){15}
//: {16}(614,379)(614,448){17}
//: {18}(#:616,450)(714,450)(714,462){19}
//: {20}(614,452)(614,511){21}
//: {22}(#:616,513)(714,513)(714,532){23}
//: {24}(614,515)(614,582){25}
//: {26}(#:616,584)(714,584)(714,601){27}
//: {28}(614,586)(614,671){29}
//: {30}(#:616,673)(714,673)(714,684){31}
//: {32}(614,675)(614,729){33}
input r6_enable;    //: /sn:0 {0}(903,280)(866,280)(866,279)(847,279){1}
input Clock_Register_File;    //: {0}(99:457,730)(556,730)(556,695){1}
//: {2}(558,693)(572,693)(572,694)(677,694){3}
//: {4}(556,691)(556,614){5}
//: {6}(558,612)(568,612)(568,611)(677,611){7}
//: {8}(556,610)(556,543){9}
//: {10}(558,541)(568,541)(568,542)(677,542){11}
//: {12}(556,539)(556,474){13}
//: {14}(558,472)(677,472){15}
//: {16}(556,470)(556,406){17}
//: {18}(558,404)(568,404)(568,403)(677,403){19}
//: {20}(556,402)(556,336){21}
//: {22}(558,334)(568,334)(568,336)(677,336){23}
//: {24}(556,332)(556,270){25}
//: {26}(558,268)(677,268){27}
//: {28}(556,266)(556,194){29}
//: {30}(558,192)(677,192){31}
//: {32}(556,190)(556,153){33}
input r3_enable;    //: /sn:0 {0}(883,487)(865,487)(865,484)(857,484){1}
input [2:0] Register_Address;    //: /sn:0 {0}(#:1166,547)(1156,547)(1156,532)(1197,532)(1197,514)(1159,514)(1159,379){1}
input r7_enable;    //: /sn:0 {0}(930,196)(882,196)(882,197)(867,197){1}
input r0_enable;    //: /sn:0 {0}(875,697)(920,697)(920,698)(930,698){1}
reg w40;    //: /sn:0 {0}(956,741)(821,741)(821,690){1}
//: {2}(821,686)(821,608){3}
//: {4}(821,604)(821,539){5}
//: {6}(821,535)(821,468){7}
//: {8}(821,464)(821,399){9}
//: {10}(821,395)(821,333){11}
//: {12}(821,329)(821,265){13}
//: {14}(821,261)(821,189){15}
//: {16}(821,185)(821,166){17}
//: {18}(819,187)(753,187){19}
//: {20}(819,263)(753,263){21}
//: {22}(819,331)(753,331){23}
//: {24}(819,397)(809,397)(809,398)(753,398){25}
//: {26}(819,466)(809,466)(809,467)(753,467){27}
//: {28}(819,537)(753,537){29}
//: {30}(819,606)(753,606){31}
//: {32}(819,688)(809,688)(809,689)(753,689){33}
wire w6;    //: /sn:0 {0}(841,484)(795,484)(50:795,477)(753,477){1}
wire [7:0] w7;    //: /sn:0 {0}(#:714,414)(714,434)(984,434){1}
//: {2}(988,434)(1041,434)(1041,352)(1143,352){3}
//: {4}(986,432)(986,409){5}
wire w4;    //: /sn:0 {0}(831,342)(784,342)(784,341)(753,341){1}
wire [7:0] w25;    //: /sn:0 {0}(#:714,203)(714,228)(1011,228){1}
//: {2}(1015,228)(#:1094,228)(1094,332)(1143,332){3}
//: {4}(1013,226)(#:1013,222)(1015,222)(1015,151){5}
wire w3;    //: /sn:0 {0}(753,197)(851,197){1}
wire [7:0] w0;    //: /sn:0 {0}(#:714,347)(714,361)(909,361)(909,345)(985,345){1}
//: {2}(989,345)(1143,345){3}
//: {4}(987,343)(987,321){5}
wire [7:0] w20;    //: /sn:0 {0}(#:714,279)(714,295)(997,295){1}
//: {2}(1001,295)(#:1082,295)(1082,339)(1143,339){3}
//: {4}(999,293)(999,273){5}
wire [7:0] w30;    //: /sn:0 {0}(#:714,622)(714,633)(987,633){1}
//: {2}(991,633)(1077,633)(1077,372)(1143,372){3}
//: {4}(989,631)(989,595){5}
wire [7:0] w10;    //: /sn:0 {0}(#:714,483)(714,492)(978,492){1}
//: {2}(982,492)(1051,492)(1051,359)(1143,359){3}
//: {4}(980,490)(#:980,480)(983,480)(983,466){5}
wire w1;    //: /sn:0 {0}(831,279)(790,279)(790,273)(753,273){1}
wire w8;    //: /sn:0 {0}(838,553)(801,553)(801,547)(753,547){1}
wire [7:0] w35;    //: /sn:0 {0}(#:714,705)(714,717)(1026,717){1}
//: {2}(1030,717)(1108,717)(1108,379)(1143,379){3}
//: {4}(1028,715)(1028,686){5}
wire w11;    //: /sn:0 {0}(859,697)(797,697)(797,699)(753,699){1}
wire [7:0] w15;    //: /sn:0 {0}(#:714,553)(714,561)(979,561){1}
//: {2}(983,561)(1061,561)(1061,365)(1143,365){3}
//: {4}(981,559)(#:981,549)(983,549)(983,532){5}
wire w5;    //: /sn:0 {0}(833,418)(805,418)(50:805,408)(753,408){1}
wire w9;    //: /sn:0 {0}(832,623)(788,623)(50:788,616)(753,616){1}
//: enddecls

  //: OUT g44 (register_file_output) @(1210,432) /sn:0 /w:[ 1 ]
  _GGREG8 #(10, 10, 20) g4 (.Q(w20), .D(register_input), .EN(w1), .CLR(w40), .CK(Clock_Register_File));   //: @(714,268) /sn:0 /w:[ 0 7 1 21 27 ]
  //: SWITCH g8 (w40) @(974,741) /sn:0 /R:2 /w:[ 0 ] /st:1 /dn:1
  _GGNBUF #(2) g47 (.I(r0_enable), .Z(w11));   //: @(869,697) /sn:0 /R:2 /w:[ 0 0 ]
  _GGREG8 #(10, 10, 20) g3 (.Q(w15), .D(register_input), .EN(w8), .CLR(w40), .CK(Clock_Register_File));   //: @(714,542) /sn:0 /w:[ 0 23 1 29 11 ]
  //: joint g16 (w40) @(821, 187) /w:[ -1 16 18 15 ]
  //: IN g26 (Clock_Register_File) @(455,730) /sn:0 /w:[ 0 ]
  //: IN g17 (r7_enable) @(932,196) /sn:0 /R:2 /w:[ 0 ]
  _GGREG8 #(10, 10, 20) g2 (.Q(w10), .D(register_input), .EN(w6), .CLR(w40), .CK(Clock_Register_File));   //: @(714,472) /sn:0 /w:[ 0 19 1 27 15 ]
  //: IN g23 (r1_enable) @(892,626) /sn:0 /R:2 /w:[ 1 ]
  //: joint g30 (Clock_Register_File) @(556, 404) /w:[ 18 20 -1 17 ]
  _GGREG8 #(10, 10, 20) g1 (.Q(w7), .D(register_input), .EN(w5), .CLR(w40), .CK(Clock_Register_File));   //: @(714,403) /sn:0 /w:[ 0 15 1 25 19 ]
  //: IN g24 (r0_enable) @(932,698) /sn:0 /R:2 /w:[ 1 ]
  //: joint g39 (register_input) @(614, 450) /w:[ 18 17 -1 20 ]
  //: LED g60 (w7) @(986,402) /sn:0 /w:[ 5 ] /type:1
  //: joint g29 (Clock_Register_File) @(556, 472) /w:[ 14 16 -1 13 ]
  _GGNBUF #(2) g51 (.I(r1_enable), .Z(w9));   //: @(842,623) /sn:0 /R:2 /w:[ 0 0 ]
  //: IN g18 (r6_enable) @(905,280) /sn:0 /R:2 /w:[ 0 ]
  //: joint g65 (w15) @(981, 561) /w:[ 2 4 1 -1 ]
  //: LED g25 (w25) @(1015,144) /sn:0 /w:[ 5 ] /type:1
  //: joint g10 (w40) @(821, 606) /w:[ -1 4 30 3 ]
  //: LED g64 (w15) @(983,525) /sn:0 /w:[ 5 ] /type:1
  _GGNBUF #(2) g49 (.I(r3_enable), .Z(w6));   //: @(851,484) /sn:0 /R:2 /w:[ 1 0 ]
  _GGNBUF #(2) g50 (.I(r2_enable), .Z(w8));   //: @(848,553) /sn:0 /R:2 /w:[ 0 0 ]
  _GGREG8 #(10, 10, 20) g6 (.Q(w30), .D(register_input), .EN(w9), .CLR(w40), .CK(Clock_Register_File));   //: @(714,611) /sn:0 /w:[ 0 27 1 31 7 ]
  //: LED g68 (w35) @(1028,679) /sn:0 /w:[ 5 ] /type:1
  //: LED g58 (w0) @(987,314) /sn:0 /w:[ 5 ] /type:1
  //: LED g56 (w20) @(999,266) /sn:0 /w:[ 5 ] /type:1
  _GGREG8 #(10, 10, 20) g7 (.Q(w35), .D(register_input), .EN(w11), .CLR(w40), .CK(Clock_Register_File));   //: @(714,694) /sn:0 /w:[ 0 31 1 33 3 ]
  //: joint g9 (w40) @(821, 688) /w:[ -1 2 32 1 ]
  //: joint g35 (register_input) @(614, 92) /w:[ 2 -1 1 4 ]
  //: joint g59 (w0) @(987, 345) /w:[ 2 4 1 -1 ]
  //: IN g22 (r2_enable) @(882,553) /sn:0 /R:2 /w:[ 1 ]
  //: joint g31 (Clock_Register_File) @(556, 334) /w:[ 22 24 -1 21 ]
  //: joint g67 (w30) @(989, 633) /w:[ 2 4 1 -1 ]
  //: joint g54 (Clock_Register_File) @(556, 693) /w:[ 2 4 -1 1 ]
  _GGMUX8x8 #(20, 20) g45 (.I0(w35), .I1(w30), .I2(w15), .I3(w10), .I4(w7), .I5(w0), .I6(w20), .I7(w25), .S(Register_Address), .Z(register_file_output));   //: @(1159,356) /sn:0 /R:1 /w:[ 3 3 3 3 3 3 3 3 1 0 ] /ss:0 /do:0
  //: joint g33 (Clock_Register_File) @(556, 192) /w:[ 30 32 -1 29 ]
  //: joint g36 (register_input) @(614, 244) /w:[ 6 5 -1 8 ]
  //: joint g41 (register_input) @(614, 584) /w:[ 26 25 -1 28 ]
  //: joint g69 (w35) @(1028, 717) /w:[ 2 4 1 -1 ]
  _GGNBUF #(2) g52 (.I(r6_enable), .Z(w1));   //: @(841,279) /sn:0 /R:2 /w:[ 1 0 ]
  //: joint g40 (register_input) @(614, 513) /w:[ 22 21 -1 24 ]
  //: joint g42 (register_input) @(614, 673) /w:[ 30 29 -1 32 ]
  //: LED g66 (w30) @(989,588) /sn:0 /w:[ 5 ] /type:1
  //: joint g12 (w40) @(821, 466) /w:[ -1 8 26 7 ]
  //: joint g57 (w20) @(999, 295) /w:[ 2 4 1 -1 ]
  //: IN g46 (Register_Address) @(1168,547) /sn:0 /R:2 /w:[ 0 ]
  //: joint g28 (Clock_Register_File) @(556, 541) /w:[ 10 12 -1 9 ]
  //: IN g34 (register_input) @(595,92) /sn:0 /w:[ 0 ]
  _GGREG8 #(10, 10, 20) g5 (.Q(w25), .D(register_input), .EN(w3), .CLR(w40), .CK(Clock_Register_File));   //: @(714,192) /sn:0 /w:[ 0 3 0 19 31 ]
  //: joint g11 (w40) @(821, 537) /w:[ -1 6 28 5 ]
  //: joint g14 (w40) @(821, 331) /w:[ -1 12 22 11 ]
  //: joint g61 (w7) @(986, 434) /w:[ 2 4 1 -1 ]
  //: IN g19 (r5_enable) @(890,341) /sn:0 /R:2 /w:[ 1 ]
  //: IN g21 (r3_enable) @(885,487) /sn:0 /R:2 /w:[ 0 ]
  //: IN g20 (r4_enable) @(903,419) /sn:0 /R:2 /w:[ 1 ]
  //: joint g32 (Clock_Register_File) @(556, 268) /w:[ 26 28 -1 25 ]
  //: joint g63 (w10) @(980, 492) /w:[ 2 4 1 -1 ]
  _GGNBUF #(2) g43 (.I(r7_enable), .Z(w3));   //: @(861,197) /sn:0 /R:2 /w:[ 1 1 ]
  _GGREG8 #(10, 10, 20) g0 (.Q(w0), .D(register_input), .EN(w4), .CLR(w40), .CK(Clock_Register_File));   //: @(714,336) /sn:0 /w:[ 0 11 1 23 23 ]
  //: joint g15 (w40) @(821, 263) /w:[ -1 14 20 13 ]
  //: joint g38 (register_input) @(614, 377) /w:[ 14 13 -1 16 ]
  _GGNBUF #(2) g48 (.I(r4_enable), .Z(w5));   //: @(843,418) /sn:0 /R:2 /w:[ 0 0 ]
  //: joint g27 (Clock_Register_File) @(556, 612) /w:[ 6 8 -1 5 ]
  //: LED g62 (w10) @(983,459) /sn:0 /w:[ 5 ] /type:1
  //: joint g37 (register_input) @(614, 303) /w:[ 10 9 -1 12 ]
  //: joint g55 (w25) @(1013, 228) /w:[ 2 4 1 -1 ]
  _GGNBUF #(2) g53 (.I(r5_enable), .Z(w4));   //: @(841,342) /sn:0 /R:2 /w:[ 0 0 ]
  //: joint g13 (w40) @(821, 397) /w:[ -1 10 24 9 ]

endmodule
//: /netlistEnd

//: /netlistBegin ram_write
module ram_write(address_to_write, write_enable, value_wrtite);
//: interface  /sz:(261, 80) /bd:[ Li0>read_addressPC[7:0](16/80) Li1>address_to_write[7:0](32/80) Li2>value_wrtite[7:0](48/80) Li3>write_enable(64/80) Ro0<w6[7:0](16/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
reg w25;    //: /sn:0 {0}(509,276)(509,281){1}
//: {2}(507,283)(497,283)(497,264){3}
//: {4}(499,262)(694,262){5}
//: {6}(497,260)(497,175){7}
//: {8}(509,285)(509,293){9}
input [7:0] address_to_write;    //: {0}(#:394,194)(99:394,235)(310,235)(310,318)(491,318){1}
reg w0;    //: /sn:0 {0}(439,525)(439,582)(468,582)(468,597){1}
input write_enable;    //: {0}(312,520)(419,520)(50:419,517)(434,517){1}
reg w2;    //: /sn:0 {0}(578,466)(578,362)(516,362)(516,343){1}
input [7:0] value_wrtite;    //: {0}(#:936,262)(50:872,262)(872,261)(862,261){1}
//: {2}(860,259)(#:860,186){3}
//: {4}(860,263)(860,326)(746,326){5}
wire w29;    //: /sn:0 {0}(439,509)(439,461)(414,461)(414,444)(434,444)(434,358)(502,358)(502,343){1}
wire w24;    //: /sn:0 {0}(710,262)(723,262)(723,341)(738,341)(738,331){1}
wire [7:0] w1;    //: /sn:0 {0}(#:526,316)(557,316)(557,326)(#:730,326){1}
//: enddecls

  _GGBUFIF8 #(4, 6) g8 (.Z(w1), .I(value_wrtite), .E(w24));   //: @(740,326) /sn:0 /R:2 /w:[ 1 5 1 ]
  _GGBUFIF #(4, 6) g4 (.Z(w29), .I(w0), .E(write_enable));   //: @(439,519) /sn:0 /R:1 /w:[ 0 0 1 ]
  //: joint g16 (w25) @(497, 262) /w:[ 4 6 -1 3 ]
  //: SWITCH g3 (w0) @(468,611) /sn:0 /R:1 /w:[ 1 ] /st:0 /dn:1
  _GGRAM8x8 #(10, 60, 70, 10, 10, 10) g26 (.A(address_to_write), .D(w1), .WE(w25), .OE(w2), .CS(w29));   //: @(509,317) /w:[ 1 0 9 1 1 ]
  //: IN g2 (address_to_write) @(394,192) /sn:0 /R:3 /w:[ 0 ]
  //: joint g1 (value_wrtite) @(860, 261) /w:[ 1 2 -1 4 ]
  //: joint g12 (w25) @(509, 283) /w:[ -1 1 2 8 ]
  //: SWITCH g11 (w2) @(578,480) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:1
  //: SWITCH g14 (w25) @(497,162) /sn:0 /R:3 /w:[ 7 ] /st:0 /dn:1
  //: IN g5 (write_enable) @(310,520) /sn:0 /w:[ 0 ]
  _GGNBUF #(2) g19 (.I(w25), .Z(w24));   //: @(700,262) /sn:0 /w:[ 5 0 ]
  //: LED g20 (value_wrtite) @(860,179) /sn:0 /w:[ 3 ] /type:1
  //: IN g0 (value_wrtite) @(938,262) /sn:0 /R:2 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin memory_read
module memory_read(w6, read_addressPC);
//: interface  /sz:(249, 40) /bd:[ Li0>read_addressPC[7:0](16/40) Ro0<w6[7:0](16/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [7:0] w6;    //: /sn:0 {0}(#:632,351)(584,351)(584,333){1}
//: {2}(584,329)(#:584,324){3}
//: {4}(582,331)(572,331)(572,287)(#:558,287)(558,227)(#:480,227){5}
reg w25;    //: /sn:0 {0}(295,101)(295,106){1}
//: {2}(293,108)(283,108)(283,0){3}
//: {4}(295,110)(295,118){5}
reg w0;    //: /sn:0 {0}(175,127)(175,114)(178,114)(178,99){1}
reg [7:0] w3;    //: /sn:0 {0}(161,167)(93,167)(#:93,203){1}
reg w29;    //: /sn:0 {0}(220,269)(220,183)(288,183)(288,168){1}
input [7:0] read_addressPC;    //: /sn:0 {0}(161,135)(122,135)(#:122,41)(#:130,41){1}
reg w2;    //: /sn:0 {0}(364,291)(364,211){1}
//: {2}(366,209)(393,209){3}
//: {4}(364,207)(364,187)(302,187)(302,168){5}
wire w7;    //: /sn:0 {0}(175,175)(175,194)(172,194)(172,209){1}
wire [7:0] w4;    //: /sn:0 {0}(#:190,151)(249,151)(249,143)(#:277,143){1}
wire [7:0] w1;    //: /sn:0 {0}(464,227)(432,227)(#:432,151)(343,151)(343,141)(#:312,141){1}
wire w28;    //: /sn:0 {0}(409,209)(472,209)(472,222){1}
//: enddecls

  //: OUT g4 (w6) @(629,351) /sn:0 /w:[ 0 ]
  //: DIP g3 (w3) @(93,214) /sn:0 /R:2 /w:[ 1 ] /st:8 /dn:1
  _GGRAM8x8 #(10, 60, 70, 10, 10, 10) g26 (.A(w4), .D(w1), .WE(w25), .OE(w2), .CS(w29));   //: @(295,142) /w:[ 1 1 5 5 1 ]
  _GGADD8 #(68, 70, 62, 64) g2 (.A(w3), .B(read_addressPC), .S(w4), .CI(w0), .CO(w7));   //: @(177,151) /sn:0 /R:1 /w:[ 0 0 0 0 0 ]
  //: SWITCH g24 (w29) @(220,283) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: IN g1 (read_addressPC) @(132,41) /sn:0 /R:2 /w:[ 1 ]
  //: joint g25 (w2) @(364, 209) /w:[ 2 4 -1 1 ]
  //: LED g6 (w7) @(172,216) /sn:0 /R:2 /w:[ 1 ] /type:0
  _GGNBUF #(2) g22 (.I(w2), .Z(w28));   //: @(399,209) /sn:0 /w:[ 3 0 ]
  //: joint g12 (w25) @(295, 108) /w:[ -1 1 2 4 ]
  //: SWITCH g5 (w0) @(178,86) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: SWITCH g11 (w2) @(364,305) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g14 (w25) @(283,-13) /sn:0 /R:3 /w:[ 3 ] /st:1 /dn:1
  _GGBUFIF8 #(4, 6) g21 (.Z(w6), .I(w1), .E(w28));   //: @(470,227) /sn:0 /w:[ 5 0 1 ]
  //: joint g0 (w6) @(584, 331) /w:[ -1 2 4 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin program_counter
module program_counter(PC_out, PC_offset, Program_counter_clock, offset_enable, PC_Clear);
//: interface  /sz:(357, 80) /bd:[ Li0>Program_counter_clock(64/80) Li1>PC_Clear(44/80) Li2>PC_offset[7:0](27/80) Li3>offset_enable(8/80) Ro0<PC_out[7:0](23/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input PC_Clear;    //: /sn:0 {0}(568,165)(568,205){1}
reg w0;    //: /sn:0 {0}(547,282)(578,282)(578,308){1}
input offset_enable;    //: /sn:0 {0}(749,346)(680,346)(680,362)(665,362){1}
reg w1;    //: /sn:0 {0}(735,528)(781,528)(781,525)(796,525){1}
input Program_counter_clock;    //: /sn:0 {0}(471,277)(423,277)(423,380){1}
output [7:0] PC_out;    //: {0}(#:508,288)(508,483)(497,483)(497,493){1}
//: {2}(499,495)(695,495)(#:695,514){3}
//: {4}(495,495)(436,495){5}
//: {6}(434,493)(434,476)(440,476)(#:50:440,457){7}
//: {8}(432,495)(394,495)(394,448){9}
reg [7:0] w5;    //: /sn:0 {0}(#:725,265)(725,315)(762,315)(762,330){1}
input [7:0] PC_offset;    //: {0}(782,330)(782,282)(#:-99:840,282){1}
wire [7:0] w6;    //: /sn:0 {0}(727,514)(727,374)(#:772,374)(#:772,359){1}
wire [7:0] w7;    //: /sn:0 {0}(508,267)(508,257)(523,257)(523,553)(711,553)(#:711,543){1}
wire w2;    //: /sn:0 {0}(568,221)(568,237)(581,237)(581,272)(547,272){1}
wire w9;    //: /sn:0 {0}(614,523)(672,523)(672,528)(687,528){1}
//: enddecls

  //: OUT g8 (PC_out) @(440,460) /sn:0 /R:1 /w:[ 7 ]
  //: LED g4 (w9) @(607,523) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: SWITCH g3 (w1) @(814,525) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  _GGMUX2x8 #(8, 8) g2 (.I0(w5), .I1(PC_offset), .S(offset_enable), .Z(w6));   //: @(772,346) /sn:0 /w:[ 1 0 0 1 ] /ss:0 /do:0
  _GGADD8 #(68, 70, 62, 64) g1 (.A(PC_out), .B(w6), .S(w7), .CI(w1), .CO(w9));   //: @(711,530) /sn:0 /w:[ 3 0 1 0 1 ]
  //: SWITCH g10 (w0) @(578,322) /sn:0 /R:1 /w:[ 1 ] /st:0 /dn:1
  //: IN g6 (PC_offset) @(842,282) /sn:0 /R:2 /w:[ 1 ]
  //: IN g7 (Program_counter_clock) @(423,382) /sn:0 /R:1 /w:[ 1 ]
  //: joint g9 (PC_out) @(434, 495) /w:[ 5 6 8 -1 ]
  //: IN g12 (offset_enable) @(663,362) /sn:0 /w:[ 1 ]
  //: LED g14 (PC_out) @(394,441) /sn:0 /w:[ 9 ] /type:1
  //: IN g11 (PC_Clear) @(568,163) /sn:0 /R:3 /w:[ 0 ]
  //: DIP g5 (w5) @(725,255) /sn:0 /w:[ 0 ] /st:2 /dn:1
  _GGREG8 #(10, 10, 20) g0 (.Q(PC_out), .D(w7), .EN(w0), .CLR(w2), .CK(Program_counter_clock));   //: @(508,277) /sn:0 /w:[ 0 0 0 1 0 ]
  //: joint g15 (PC_out) @(497, 495) /w:[ 2 1 4 -1 ]
  _GGNBUF #(2) g13 (.I(PC_Clear), .Z(w2));   //: @(568,211) /sn:0 /R:3 /w:[ 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin xor_gate
module xor_gate(xor_gate_output, xor_gate_input_2, xor_gate_input_1, xor_enable);
//: interface  /sz:(255, 64) /bd:[ Li0>xor_enable(48/64) Li1>xor_gate_input_2[7:0](32/64) Li2>xor_gate_input_1[7:0](16/64) Ro0<xor_gate_output[7:0](16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] xor_gate_input_1;    //: /sn:0 {0}(232,134)(232,120)(#:202,120){1}
input [7:0] xor_gate_input_2;    //: /sn:0 {0}(254,216)(254,243)(#:222,243)(#:222,256)(#:207,256){1}
input xor_enable;    //: /sn:0 {0}(249,208)(77,208)(77,186){1}
//: {2}(77,182)(77,157)(247,157)(247,142)(237,142){3}
//: {4}(75,184)(62,184){5}
output [7:0] xor_gate_output;    //: {0}(#:348,178)(371,178)(96:371,179)(510,179){1}
wire [7:0] w0;    //: /sn:0 {0}(#:254,200)(254,180)(#:50:327,180){1}
wire [7:0] w1;    //: /sn:0 {0}(#:232,150)(232,175)(#:50:327,175){1}
//: enddecls

  _GGBUFIF8 #(4, 6) g4 (.Z(w1), .I(xor_gate_input_1), .E(xor_enable));   //: @(232,140) /sn:0 /R:3 /w:[ 0 0 3 ]
  //: OUT g3 (xor_gate_output) @(507,179) /sn:0 /w:[ 1 ]
  //: IN g2 (xor_gate_input_2) @(205,256) /sn:0 /w:[ 1 ]
  //: IN g1 (xor_gate_input_1) @(200,120) /sn:0 /w:[ 1 ]
  //: IN g6 (xor_enable) @(60,184) /sn:0 /w:[ 5 ]
  //: joint g7 (xor_enable) @(77, 184) /w:[ -1 2 4 1 ]
  _GGBUFIF8 #(4, 6) g5 (.Z(w0), .I(xor_gate_input_2), .E(xor_enable));   //: @(254,210) /sn:0 /R:1 /w:[ 0 0 0 ]
  _GGXOR2x8 #(8) g0 (.I0(w1), .I1(w0), .Z(xor_gate_output));   //: @(338,178) /sn:0 /w:[ 1 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin comparator
module comparator(input_2, input_1, comparator_enable, comparator_result);
//: interface  /sz:(279, 64) /bd:[ Li0>comparator_enable(48/64) Li1>input_2[7:0](32/64) Li2>input_1[7:0](16/64) Ro0<comparator_result(16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] input_1;    //: {0}(#:-80:495,277)(#:509,277)(509,295)(524,295){1}
input comparator_enable;    //: {0}(532,290)(532,278)(517,278)(517,324){1}
//: {2}(519,326)(537,326)(537,348){3}
//: {4}(98:515,326)(408,326){5}
input [7:0] input_2;    //: /sn:0 {0}(#:500,389)(#:514,389)(514,353)(529,353){1}
output comparator_result;    //: {0}(918,348)(942,348)(942,336)(50:952,336){1}
wire w6;    //: /sn:0 {0}(897,356)(778,356){1}
//: {2}(776,354)(776,289){3}
//: {4}(776,358)(776,405)(642,405){5}
wire w7;    //: /sn:0 {0}(897,361)(803,361)(803,362)(793,362){1}
//: {2}(791,360)(791,289){3}
//: {4}(791,364)(791,425)(642,425){5}
wire w4;    //: /sn:0 {0}(897,346)(746,346){1}
//: {2}(744,344)(744,289){3}
//: {4}(744,348)(744,367)(642,367){5}
wire w3;    //: /sn:0 {0}(897,341)(731,341){1}
//: {2}(729,339)(729,289){3}
//: {4}(729,343)(729,349)(642,349){5}
wire w0;    //: /sn:0 {0}(642,314)(679,314){1}
//: {2}(683,314)(697,314)(697,289){3}
//: {4}(681,316)(681,331)(897,331){5}
wire [7:0] w10;    //: /sn:0 {0}(#:545,353)(563,353)(563,307)(#:597,307){1}
wire w1;    //: /sn:0 {0}(642,332)(668,332){1}
//: {2}(672,332)(714,332)(714,289){3}
//: {4}(670,334)(670,336)(897,336){5}
wire w8;    //: /sn:0 {0}(897,366)(810,366){1}
//: {2}(808,364)(808,289){3}
//: {4}(808,368)(808,442)(642,442){5}
wire [7:0] w2;    //: /sn:0 {0}(#:618,305)(638,305)(638,313){1}
//: {2}(638,314)(638,331){3}
//: {4}(638,332)(638,348){5}
//: {6}(638,349)(638,366){7}
//: {8}(638,367)(638,385){9}
//: {10}(638,386)(638,404){11}
//: {12}(638,405)(638,424){13}
//: {14}(638,425)(638,441){15}
//: {16}(638,442)(638,450){17}
wire w5;    //: /sn:0 {0}(897,351)(773,351)(773,350)(763,350){1}
//: {2}(761,348)(761,289){3}
//: {4}(761,352)(761,386)(642,386){5}
wire [7:0] w9;    //: /sn:0 {0}(#:540,295)(552,295)(552,302)(#:597,302){1}
//: enddecls

  //: LED g8 (w4) @(744,282) /sn:0 /w:[ 3 ] /type:1
  assign w0 = w2[0]; //: TAP g4 @(636,314) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  assign w7 = w2[6]; //: TAP g16 @(636,425) /sn:0 /R:2 /w:[ 5 14 13 ] /ss:1
  //: LED g3 (w0) @(697,282) /sn:0 /w:[ 3 ] /type:1
  //: joint g26 (w7) @(791, 362) /w:[ 1 2 -1 4 ]
  //: LED g17 (w8) @(808,282) /sn:0 /w:[ 3 ] /type:1
  //: IN g2 (input_2) @(498,389) /sn:0 /w:[ 0 ]
  _GGBUFIF8 #(4, 6) g30 (.Z(w10), .I(input_2), .E(comparator_enable));   //: @(535,353) /sn:0 /w:[ 0 1 3 ]
  //: joint g23 (w4) @(744, 346) /w:[ 1 2 -1 4 ]
  //: joint g24 (w5) @(761, 350) /w:[ 1 2 -1 4 ]
  //: IN g1 (input_1) @(493,277) /sn:0 /w:[ 0 ]
  _GGBUFIF8 #(4, 6) g29 (.Z(w9), .I(input_1), .E(comparator_enable));   //: @(530,295) /sn:0 /w:[ 0 1 0 ]
  assign w8 = w2[7]; //: TAP g18 @(636,442) /sn:0 /R:2 /w:[ 5 16 15 ] /ss:1
  //: joint g25 (w6) @(776, 356) /w:[ 1 2 -1 4 ]
  //: LED g10 (w6) @(776,282) /sn:0 /w:[ 3 ] /type:1
  assign w1 = w2[1]; //: TAP g6 @(636,332) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: LED g9 (w5) @(761,282) /sn:0 /w:[ 3 ] /type:1
  //: LED g7 (w3) @(729,282) /sn:0 /w:[ 3 ] /type:1
  //: IN g31 (comparator_enable) @(406,326) /sn:0 /w:[ 5 ]
  //: joint g22 (w3) @(729, 341) /w:[ 1 2 -1 4 ]
  assign w3 = w2[2]; //: TAP g12 @(636,349) /sn:0 /R:2 /w:[ 5 6 5 ] /ss:1
  //: OUT g28 (comparator_result) @(949,336) /sn:0 /w:[ 1 ]
  assign w5 = w2[4]; //: TAP g14 @(636,386) /sn:0 /R:2 /w:[ 5 10 9 ] /ss:1
  //: LED g11 (w7) @(791,282) /sn:0 /w:[ 3 ] /type:1
  //: LED g5 (w1) @(714,282) /sn:0 /w:[ 3 ] /type:1
  //: joint g21 (w1) @(670, 332) /w:[ 2 -1 1 4 ]
  _GGOR8 #(18) g19 (.I0(w0), .I1(w1), .I2(w3), .I3(w4), .I4(w5), .I5(w6), .I6(w7), .I7(w8), .Z(comparator_result));   //: @(908,348) /sn:0 /w:[ 5 5 0 0 0 0 0 0 0 ]
  //: joint g32 (comparator_enable) @(517, 326) /w:[ 2 1 4 -1 ]
  //: joint g20 (w0) @(681, 314) /w:[ 2 -1 1 4 ]
  assign w6 = w2[5]; //: TAP g15 @(636,405) /sn:0 /R:2 /w:[ 5 12 11 ] /ss:1
  _GGXOR2x8 #(8) g0 (.I0(w9), .I1(w10), .Z(w2));   //: @(608,305) /sn:0 /w:[ 1 1 0 ]
  //: joint g27 (w8) @(808, 366) /w:[ 1 2 -1 4 ]
  assign w4 = w2[3]; //: TAP g13 @(636,367) /sn:0 /R:2 /w:[ 5 8 7 ] /ss:1

endmodule
//: /netlistEnd

